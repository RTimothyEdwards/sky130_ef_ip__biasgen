magic
tech sky130A
magscale 1 2
timestamp 1747752771
<< locali >>
rect 1986 -3003 2210 -2709
rect 2470 -2752 2520 -2709
rect 2470 -2945 2480 -2752
rect 2514 -2945 2520 -2752
rect 2470 -3003 2520 -2945
<< viali >>
rect 2480 -2945 2514 -2752
<< metal1 >>
rect 2062 244 2641 302
rect 2062 234 2122 244
rect 2063 166 2122 234
rect 2588 166 2641 244
rect 2063 154 2641 166
rect 2063 -1889 2115 154
rect 2150 -1478 2214 8
rect 2326 -565 2378 92
rect 2482 14 2641 154
rect 2470 -582 2641 14
rect 2326 -757 2378 -751
rect 2325 -1463 2377 -802
rect 2325 -1654 2377 -1648
rect 2330 -1707 2378 -1700
rect 2059 -2406 2111 -1889
rect 2059 -2548 2111 -2542
rect 2144 -3439 2208 -1772
rect 2144 -3697 2208 -3671
rect 2330 -3132 2384 -1707
rect 2480 -2360 2544 -887
rect 2589 -1889 2641 -582
rect 2593 -2406 2645 -1889
rect 2593 -2551 2645 -2542
rect 2470 -2731 2540 -2709
rect 2470 -3003 2540 -2969
rect 2330 -3697 2384 -3364
<< via1 >>
rect 2122 166 2588 244
rect 2326 -751 2378 -565
rect 2325 -1648 2377 -1463
rect 2059 -2542 2111 -2406
rect 2144 -3671 2208 -3439
rect 2593 -2542 2645 -2406
rect 2470 -2752 2540 -2731
rect 2470 -2945 2480 -2752
rect 2480 -2945 2514 -2752
rect 2514 -2945 2540 -2752
rect 2470 -2969 2540 -2945
rect 2330 -3364 2384 -3132
<< metal2 >>
rect 1986 244 2714 338
rect 1986 166 2122 244
rect 2588 166 2714 244
rect 1986 104 2714 166
rect 2326 -565 2378 -558
rect 1986 -751 2326 -608
rect 2378 -751 2714 -608
rect 1986 -842 2714 -751
rect 2325 -1463 2377 -1457
rect 1986 -1648 2325 -1507
rect 2377 -1648 2714 -1507
rect 1986 -1741 2714 -1648
rect 1986 -2406 2714 -2400
rect 1986 -2542 2059 -2406
rect 2111 -2542 2593 -2406
rect 2645 -2542 2714 -2406
rect 1986 -2634 2714 -2542
rect 1986 -2969 2470 -2731
rect 2540 -2969 2714 -2731
rect 2324 -3364 2330 -3132
rect 2384 -3364 2390 -3132
rect 2138 -3671 2144 -3439
rect 2208 -3671 2214 -3439
use sky130_fd_pr__diode_pw2nd_05v5_FT76RK  sky130_fd_pr__diode_pw2nd_05v5_FT76RK_0 paramcells
timestamp 1713888873
transform 1 0 2357 0 1 -2856
box -183 -183 183 183
use sky130_fd_pr__pfet_g5v0d10v5_G8LMTE  sky130_fd_pr__pfet_g5v0d10v5_G8LMTE_0 paramcells
timestamp 1747745073
transform 1 0 2352 0 1 -2073
box -362 -550 362 543
use sky130_fd_pr__pfet_g5v0d10v5_H75TTF  sky130_fd_pr__pfet_g5v0d10v5_H75TTF_0 paramcells
timestamp 1747745073
transform 1 0 2352 0 1 -281
box -362 -543 362 547
use sky130_fd_pr__pfet_g5v0d10v5_G8LMTE  XM13
timestamp 1747745073
transform 1 0 2352 0 1 -1177
box -362 -550 362 543
<< labels >>
flabel metal1 2480 -1662 2544 -1600 0 FreeSans 560 90 0 0 vcasc
port 7 nsew
flabel metal2 1990 104 2122 338 0 FreeSans 560 0 0 0 avdd
port 0 nsew
flabel metal2 2540 -2969 2710 -2731 0 FreeSans 560 0 0 0 avss
port 1 nsew
flabel metal1 2330 -3697 2384 -3526 0 FreeSans 560 90 0 0 enb
port 4 nsew
flabel metal1 2144 -3388 2208 -3218 0 FreeSans 560 90 0 0 itail
port 5 nsew
flabel metal2 1990 -1741 2326 -1507 0 FreeSans 560 0 0 0 pcasc
port 3 nsew
flabel metal2 2378 -842 2710 -608 0 FreeSans 560 0 0 0 pbias
port 8 nsew
<< end >>
