magic
tech sky130A
magscale 1 2
timestamp 1747745286
<< locali >>
rect 3392 114 3448 408
rect 3742 114 3926 408
rect 3392 92 3926 114
rect 3448 20 3742 92
<< metal1 >>
rect 3724 777 3788 785
rect 3568 521 3622 527
rect 3300 30 3352 40
rect 3352 -106 3353 26
rect 3300 -112 3353 -106
rect 3301 -1916 3353 -112
rect 3392 -1611 3456 -119
rect 3568 -784 3622 333
rect 3724 -726 3788 589
rect 3834 32 3886 40
rect 3834 30 3887 32
rect 3886 -106 3887 30
rect 3834 -112 3887 -106
rect 3568 -1667 3620 -938
rect 3301 -2632 3456 -1916
rect 3568 -2584 3620 -1863
rect 3726 -2502 3790 -1019
rect 3568 -2586 3616 -2584
rect 3835 -2632 3887 -112
rect 3301 -2690 3887 -2632
rect 3300 -2704 3890 -2690
rect 3300 -2782 3358 -2704
rect 3832 -2782 3890 -2704
rect 3300 -2796 3890 -2782
<< via1 >>
rect 3724 589 3788 777
rect 3568 333 3622 521
rect 3300 -106 3352 30
rect 3834 -106 3886 30
rect 3568 -1863 3620 -1667
rect 3358 -2782 3832 -2704
<< metal2 >>
rect 3718 589 3724 777
rect 3788 589 3794 777
rect 3560 333 3568 521
rect 3622 333 3631 521
rect 3258 30 3926 124
rect 3258 -106 3300 30
rect 3352 -106 3834 30
rect 3886 -106 3926 30
rect 3258 -114 3926 -106
rect 3258 -1667 3926 -1643
rect 3258 -1863 3568 -1667
rect 3620 -1863 3926 -1667
rect 3258 -1881 3926 -1863
rect 3258 -2704 3926 -2622
rect 3258 -2782 3358 -2704
rect 3832 -2782 3926 -2704
rect 3258 -2860 3926 -2782
use sky130_fd_pr__diode_pw2nd_05v5_FT76RK  sky130_fd_pr__diode_pw2nd_05v5_FT76RK_0 paramcells
timestamp 1713888873
transform 1 0 3595 0 1 261
box -183 -183 183 183
use sky130_fd_pr__nfet_05v0_nvt_QRKT8A  XM6 paramcells
timestamp 1747745286
transform 1 0 3594 0 1 -1316
box -332 -513 332 513
use sky130_fd_pr__nfet_g5v0d10v5_ZMKT8B  XM7 paramcells
timestamp 1747745286
transform 1 0 3594 0 1 -420
box -332 -513 332 513
use sky130_fd_pr__nfet_g5v0d10v5_C3WBNC  XM12 paramcells
timestamp 1747745286
transform 1 0 3594 0 1 -2212
box -332 -513 332 513
<< labels >>
flabel metal1 3392 -612 3456 -550 0 FreeSans 560 90 0 0 vcasc
port 5 nsew
flabel metal2 3258 -2860 3358 -2622 0 FreeSans 560 90 0 0 avss
port 1 nsew
flabel metal2 3262 -1881 3568 -1643 0 FreeSans 560 0 0 0 nbias
port 4 nsew
flabel metal1 3568 154 3622 208 0 FreeSans 560 0 0 0 ena
port 3 nsew
flabel metal1 3724 440 3788 542 0 FreeSans 560 90 0 0 itail
port 2 nsew
<< end >>
