magic
tech sky130A
magscale 1 2
timestamp 1719970077
<< error_s >>
rect 45076 7047 45976 7947
<< dnwell >>
rect 5006 301 45976 8153
<< nwell >>
rect 4897 7947 45976 8262
rect 4897 507 5212 7947
rect 4897 192 45976 507
<< pwell >>
rect 19789 766 19859 1198
rect 35342 507 35430 529
<< mvpsubdiff >>
rect 4777 8352 4837 8386
rect 45787 8352 45910 8386
rect 4777 8326 4811 8352
rect 1075 7702 1135 7736
rect 4170 7702 4230 7736
rect 1075 7676 1109 7702
rect 1075 682 1109 708
rect 4196 7676 4230 7702
rect 4196 682 4230 708
rect 1075 648 1135 682
rect 4170 648 4230 682
rect 4777 80 4811 106
rect 4777 46 4837 80
rect 45777 46 45910 80
<< mvnsubdiff >>
rect 4963 8176 45910 8196
rect 4963 8142 5043 8176
rect 45787 8142 45910 8176
rect 4963 8122 45910 8142
rect 4963 8116 5037 8122
rect 4963 338 4983 8116
rect 5017 338 5037 8116
rect 4963 332 5037 338
rect 4963 312 45910 332
rect 4963 278 5043 312
rect 45777 278 45910 312
rect 4963 258 45910 278
<< mvpsubdiffcont >>
rect 4837 8352 45787 8386
rect 1135 7702 4170 7736
rect 1075 708 1109 7676
rect 4196 708 4230 7676
rect 1135 648 4170 682
rect 4777 106 4811 8326
rect 4837 46 45777 80
<< mvnsubdiffcont >>
rect 5043 8142 45787 8176
rect 4983 338 5017 8116
rect 5043 278 45777 312
<< locali >>
rect 4777 8352 4837 8386
rect 45787 8352 45910 8386
rect 4777 8326 45910 8352
rect 1072 7736 4777 7837
rect 1072 7702 1135 7736
rect 4170 7713 4777 7736
rect 4170 7702 4341 7713
rect 1072 7676 1209 7702
rect 1072 708 1075 7676
rect 1109 708 1209 7676
rect 4196 7676 4341 7702
rect 3464 7097 3511 7163
rect 1707 6273 1873 6285
rect 1707 6164 1720 6273
rect 1857 6164 1873 6273
rect 1707 6151 1873 6164
rect 1707 4645 1873 4657
rect 1707 4536 1720 4645
rect 1857 4536 1873 4645
rect 1707 4523 1873 4536
rect 3464 3841 3511 3907
rect 1707 3017 1873 3029
rect 1707 2908 1720 3017
rect 1857 2908 1873 3017
rect 1707 2895 1873 2908
rect 1707 1389 1873 1401
rect 1707 1280 1720 1389
rect 1857 1280 1873 1389
rect 1707 1267 1873 1280
rect 1072 682 1209 708
rect 4230 708 4341 7676
rect 4196 682 4341 708
rect 4811 8253 45910 8326
rect 4811 2306 4879 8253
rect 1072 648 1135 682
rect 4170 648 4777 682
rect 1072 558 4777 648
rect 4852 224 4879 2306
rect 4983 8142 5043 8176
rect 45787 8142 45902 8176
rect 4983 8116 45902 8142
rect 5017 7957 45902 8116
rect 5017 7498 5151 7957
rect 5136 7294 5151 7498
rect 5017 5883 5151 7294
rect 5017 4240 5019 5883
rect 5128 4240 5151 5883
rect 5906 5647 6200 5658
rect 5906 5570 5917 5647
rect 6187 5570 6200 5647
rect 5906 5561 6200 5570
rect 5017 491 5151 4240
rect 5017 338 45902 491
rect 4983 312 45902 338
rect 4983 278 5043 312
rect 45777 278 45902 312
rect 4811 192 4879 224
rect 4811 106 45910 192
rect 4777 105 45910 106
rect 4777 61 4804 105
rect 4777 46 4837 61
rect 45777 46 45910 105
<< viali >>
rect 3782 7073 3848 7300
rect 3398 6825 3464 7052
rect 1720 6164 1857 6273
rect 3398 5197 3464 5424
rect 1720 4536 1857 4645
rect 3782 3817 3848 4044
rect 1720 2908 1857 3017
rect 3398 1941 3464 2168
rect 1720 1280 1857 1389
rect 4803 224 4811 2306
rect 4811 224 4852 2306
rect 4999 7294 5017 7498
rect 5017 7294 5136 7498
rect 5019 4240 5128 5883
rect 5917 5570 6187 5647
rect 4804 80 45777 105
rect 4804 61 4837 80
rect 4837 61 45777 80
<< metal1 >>
rect 1371 7535 3964 7554
rect 1371 7409 1559 7535
rect 2043 7409 3964 7535
rect 1371 7391 3964 7409
rect 4982 7498 5151 7512
rect 3775 7300 3856 7317
rect 3775 7073 3782 7300
rect 3848 7175 3856 7300
rect 4370 7175 4376 7344
rect 3848 7112 4376 7175
rect 3848 7073 3856 7112
rect 4370 7111 4376 7112
rect 4434 7175 4440 7344
rect 4730 7175 4736 7344
rect 4434 7112 4736 7175
rect 4434 7111 4440 7112
rect 4730 7111 4736 7112
rect 4794 7111 4800 7344
rect 4982 7294 4999 7498
rect 5136 7294 5151 7498
rect 4982 7278 5151 7294
rect 3391 7052 3472 7069
rect 3775 7060 3856 7073
rect 3391 6825 3398 7052
rect 3464 6938 3472 7052
rect 4490 6938 4496 7024
rect 3464 6880 4496 6938
rect 3464 6825 3472 6880
rect 3391 6812 3472 6825
rect 4490 6791 4496 6880
rect 4554 6938 4560 7024
rect 4554 6880 4577 6938
rect 4554 6791 4560 6880
rect 1378 6717 3971 6741
rect 1378 6591 3158 6717
rect 3642 6591 3971 6717
rect 1378 6578 3971 6591
rect 1707 6273 1873 6285
rect 1707 6253 1720 6273
rect 1072 6185 1720 6253
rect 1707 6164 1720 6185
rect 1857 6164 1873 6273
rect 1707 6151 1873 6164
rect 1368 5906 3961 5921
rect 1368 5780 1560 5906
rect 2044 5780 3961 5906
rect 1368 5758 3961 5780
rect 5002 5883 5149 5901
rect 3391 5424 3472 5441
rect 3391 5197 3398 5424
rect 3464 5310 3472 5424
rect 4490 5310 4496 5495
rect 3464 5262 4496 5310
rect 4554 5310 4560 5495
rect 4554 5262 4577 5310
rect 3464 5252 4577 5262
rect 3464 5197 3472 5252
rect 3391 5184 3472 5197
rect 1376 5094 3969 5113
rect 1376 4968 3162 5094
rect 3646 4968 3969 5094
rect 1376 4950 3969 4968
rect 1707 4645 1873 4657
rect 1707 4625 1720 4645
rect 1072 4557 1720 4625
rect 1707 4536 1720 4557
rect 1857 4536 1873 4645
rect 1707 4523 1873 4536
rect 1368 4266 3961 4288
rect 1368 4140 1557 4266
rect 2041 4140 3961 4266
rect 5002 4240 5019 5883
rect 5128 4240 5149 5883
rect 5441 5459 5562 8557
rect 19859 7753 33103 7764
rect 19859 7701 19892 7753
rect 33067 7701 33103 7753
rect 19859 7689 33103 7701
rect 8071 7171 8491 7593
rect 8071 6504 8242 7171
rect 8597 7166 8833 7598
rect 8929 7166 9165 7598
rect 9261 7166 9497 7598
rect 9593 7166 9829 7598
rect 9925 7166 10161 7598
rect 10257 7166 10493 7598
rect 10589 7166 10825 7598
rect 10921 7166 11157 7598
rect 11253 7166 11489 7598
rect 11585 7166 11821 7598
rect 11917 7166 12153 7598
rect 12249 7166 12485 7598
rect 12581 7166 12817 7598
rect 12913 7166 13149 7598
rect 13245 7166 13481 7598
rect 13577 7166 13813 7598
rect 13909 7166 14145 7598
rect 14241 7166 14477 7598
rect 14573 7166 14809 7598
rect 14905 7166 15141 7598
rect 15237 7166 15473 7598
rect 15569 7166 15805 7598
rect 15901 7166 16137 7598
rect 16233 7166 16469 7598
rect 16565 7166 16801 7598
rect 16897 7166 17133 7598
rect 17229 7166 17465 7598
rect 17561 7166 17797 7598
rect 17893 7166 18129 7598
rect 18225 7166 18461 7598
rect 18557 7166 18793 7598
rect 18889 7166 19125 7598
rect 19221 7166 19457 7598
rect 6727 6333 8242 6504
rect 6727 6226 6898 6333
rect 5747 6215 6898 6226
rect 5747 6067 5761 6215
rect 6157 6067 6898 6215
rect 5747 6055 6898 6067
rect 5896 5647 8331 5658
rect 5896 5570 5917 5647
rect 6187 5570 8331 5647
rect 5896 5561 8331 5570
rect 5441 5426 6822 5459
rect 5002 4218 5149 4240
rect 5557 4356 5651 4367
rect 1368 4125 3961 4140
rect 5557 4141 5566 4356
rect 5639 4141 5651 4356
rect 6789 4184 6822 5426
rect 5557 4131 5651 4141
rect 3775 4044 3856 4061
rect 3775 3817 3782 4044
rect 3848 3921 3856 4044
rect 4610 3921 4616 4106
rect 3848 3873 4616 3921
rect 4674 3873 4680 4106
rect 3848 3864 4680 3873
rect 3848 3817 3856 3864
rect 3775 3804 3856 3817
rect 1373 3460 3966 3482
rect 1373 3334 3160 3460
rect 3644 3334 3966 3460
rect 1373 3319 3966 3334
rect 1707 3017 1873 3029
rect 1707 2997 1720 3017
rect 1072 2929 1720 2997
rect 1707 2908 1720 2929
rect 1857 2908 1873 3017
rect 1707 2895 1873 2908
rect 1371 2648 3964 2669
rect 1371 2522 1558 2648
rect 2042 2522 3964 2648
rect 1371 2506 3964 2522
rect 4777 2306 4879 2345
rect 3391 2168 3472 2185
rect 3391 1941 3398 2168
rect 3464 2054 3472 2168
rect 4490 2054 4496 2229
rect 3464 1996 4496 2054
rect 4554 2054 4560 2229
rect 4777 2181 4803 2306
rect 4554 1996 4577 2054
rect 3464 1941 3472 1996
rect 3391 1928 3472 1941
rect 1371 1832 3966 1856
rect 1371 1706 3158 1832
rect 3642 1706 3966 1832
rect 1371 1691 3966 1706
rect 1707 1389 1873 1401
rect 1707 1369 1720 1389
rect 1072 1301 1720 1369
rect 1707 1280 1720 1301
rect 1857 1280 1873 1389
rect 1707 1267 1873 1280
rect 1380 970 1560 1035
rect 2044 970 3963 1035
rect 4775 622 4803 2181
rect 4777 224 4803 622
rect 4852 2181 4879 2306
rect 4852 2161 5211 2181
rect 4852 641 5042 2161
rect 5198 641 5211 2161
rect 19541 1546 19593 7598
rect 19789 7166 20025 7598
rect 20121 7166 20357 7598
rect 20453 7166 20689 7598
rect 20785 7166 21021 7598
rect 21117 7166 21353 7598
rect 21449 7166 21685 7598
rect 21781 7166 22017 7598
rect 22113 7166 22349 7598
rect 22445 7166 22681 7598
rect 22777 7166 23013 7598
rect 23109 7166 23345 7598
rect 23441 7166 23677 7598
rect 23773 7166 24009 7598
rect 24105 7166 24341 7598
rect 24437 7166 24673 7598
rect 24769 7166 25005 7598
rect 25101 7166 25337 7598
rect 25433 7166 25669 7598
rect 25765 7166 26001 7598
rect 26097 7166 26333 7598
rect 26429 7166 26665 7598
rect 26761 7166 26997 7598
rect 27093 7166 27329 7598
rect 27425 7166 27661 7598
rect 27757 7166 27993 7598
rect 28089 7166 28325 7598
rect 28421 7166 28657 7598
rect 28753 7166 28989 7598
rect 29085 7166 29321 7598
rect 29417 7166 29653 7598
rect 29749 7166 29985 7598
rect 30081 7166 30317 7598
rect 30413 7166 30649 7598
rect 30745 7166 30981 7598
rect 31077 7166 31313 7598
rect 31409 7166 31645 7598
rect 31741 7166 31977 7598
rect 32073 7166 32309 7598
rect 32405 7166 32641 7598
rect 32737 7166 32973 7598
rect 19541 1198 19593 1308
rect 19653 1546 19705 7004
rect 19653 1296 19705 1308
rect 27923 6512 28159 6521
rect 8431 766 8667 1198
rect 8763 766 8999 1198
rect 9095 766 9331 1198
rect 9427 766 9663 1198
rect 9759 766 9995 1198
rect 10091 766 10327 1198
rect 10423 766 10659 1198
rect 10755 766 10991 1198
rect 11087 766 11323 1198
rect 11419 766 11655 1198
rect 11751 766 11987 1198
rect 12083 766 12319 1198
rect 12415 766 12651 1198
rect 12747 766 12983 1198
rect 13079 766 13315 1198
rect 13411 766 13647 1198
rect 13743 766 13979 1198
rect 14075 766 14311 1198
rect 14407 766 14643 1198
rect 14739 766 14975 1198
rect 15071 766 15307 1198
rect 15403 766 15639 1198
rect 15735 766 15971 1198
rect 16067 766 16303 1198
rect 16399 766 16635 1198
rect 16731 766 16967 1198
rect 17063 766 17299 1198
rect 17395 766 17631 1198
rect 17727 766 17963 1198
rect 18059 766 18295 1198
rect 18391 766 18627 1198
rect 18723 766 18959 1198
rect 19055 766 19291 1198
rect 19387 766 19593 1198
rect 19641 1189 19859 1198
rect 19641 776 19652 1189
rect 19748 776 19859 1189
rect 19641 766 19859 776
rect 19955 766 20191 1198
rect 20287 766 20523 1198
rect 20619 766 20855 1198
rect 20951 766 21187 1198
rect 21283 766 21519 1198
rect 21615 766 21851 1198
rect 21947 766 22183 1198
rect 22279 766 22515 1198
rect 22611 766 22847 1198
rect 22943 766 23179 1198
rect 23275 766 23511 1198
rect 23607 766 23843 1198
rect 23939 766 24175 1198
rect 24271 766 24507 1198
rect 24603 766 24839 1198
rect 24935 766 25171 1198
rect 25267 766 25503 1198
rect 25599 766 25835 1198
rect 25931 766 26167 1198
rect 26263 766 26499 1198
rect 26595 766 26831 1198
rect 26927 766 27163 1198
rect 27259 766 27495 1198
rect 27591 766 27827 1198
rect 27923 766 28159 6278
rect 33063 4062 33115 4076
rect 33063 3810 33115 3824
rect 34878 2716 35072 2800
rect 35412 2716 35606 2800
rect 35946 2716 36140 2800
rect 36480 2716 36674 2800
rect 37014 2716 37208 2800
rect 37548 2716 37742 2800
rect 38082 2716 38276 2800
rect 38616 2716 38810 2800
rect 39150 2716 39344 2800
rect 39684 2716 39878 2800
rect 40218 2716 40412 2800
rect 40752 2716 40946 2800
rect 41286 2716 41480 2800
rect 41820 2716 42014 2800
rect 42354 2716 42548 2800
rect 42888 2716 43082 2800
rect 43422 2716 43616 2800
rect 43956 2716 44150 2800
rect 44490 2716 44684 2800
rect 45024 2716 45218 2800
rect 28255 766 28491 1198
rect 28587 766 28823 1198
rect 28919 766 29155 1198
rect 29251 766 29487 1198
rect 29583 766 29819 1198
rect 29915 766 30151 1198
rect 30247 766 30483 1198
rect 30579 766 30815 1198
rect 30911 766 31147 1198
rect 31243 766 31479 1198
rect 31575 766 31811 1198
rect 31907 766 32143 1198
rect 32239 766 32475 1198
rect 32571 766 32807 1198
rect 32903 1190 33107 1198
rect 32903 776 33009 1190
rect 33096 776 33107 1190
rect 32903 766 33107 776
rect 4852 622 5211 641
rect 19541 630 19593 766
rect 4852 224 4879 622
rect 4777 124 4879 224
rect 4777 105 45900 124
rect 4777 61 4804 105
rect 45777 61 45900 105
rect 4777 46 45900 61
<< via1 >>
rect 1559 7409 2043 7535
rect 4376 7111 4434 7344
rect 4736 7111 4794 7344
rect 4999 7294 5136 7498
rect 4496 6791 4554 7024
rect 3158 6591 3642 6717
rect 2348 6449 2858 6506
rect 1560 5780 2044 5906
rect 4496 5262 4554 5495
rect 3162 4968 3646 5094
rect 2348 4821 2858 4878
rect 1557 4140 2041 4266
rect 5019 4240 5128 5883
rect 19892 7701 33067 7753
rect 5761 6067 6157 6215
rect 5566 4141 5639 4356
rect 4616 3873 4674 4106
rect 3160 3334 3644 3460
rect 2348 3193 2858 3250
rect 1558 2522 2042 2648
rect 4496 1996 4554 2229
rect 3158 1706 3642 1832
rect 2348 1565 2858 1622
rect 1560 956 2044 1070
rect 5042 641 5198 2161
rect 19541 1308 19593 1546
rect 19653 1308 19705 1546
rect 27923 6278 28159 6512
rect 19652 776 19748 1189
rect 33063 3824 33115 4062
rect 33009 776 33096 1190
<< metal2 >>
rect 33214 8636 45248 8715
rect 33214 8250 33293 8636
rect 33578 8317 33721 8549
rect 33927 8317 38469 8549
rect 38905 8539 44901 8549
rect 38905 8326 38920 8539
rect 38989 8326 39454 8539
rect 39523 8326 39988 8539
rect 40057 8326 40522 8539
rect 40591 8326 41056 8539
rect 41125 8326 41590 8539
rect 41659 8326 42124 8539
rect 42193 8326 42658 8539
rect 42727 8326 43192 8539
rect 43261 8326 43726 8539
rect 43795 8326 44260 8539
rect 44329 8326 44794 8539
rect 44863 8326 44901 8539
rect 38905 8317 44901 8326
rect 4496 8171 33293 8250
rect 45169 8242 45248 8636
rect 45302 8535 45609 8549
rect 45302 8332 45318 8535
rect 45595 8332 45609 8535
rect 45302 8317 45609 8332
rect 1548 7535 2059 7630
rect 1548 7409 1559 7535
rect 2043 7409 2059 7535
rect 1548 5906 2059 7409
rect 1548 5780 1560 5906
rect 2044 5780 2059 5906
rect 1548 4266 2059 5780
rect 1548 4140 1557 4266
rect 2041 4140 2059 4266
rect 1548 2648 2059 4140
rect 1548 2522 1558 2648
rect 2042 2522 2059 2648
rect 1548 2096 2059 2522
rect 1548 1489 1582 2096
rect 2027 1489 2059 2096
rect 1548 1070 2059 1489
rect 1548 956 1560 1070
rect 2044 956 2059 1070
rect 1548 820 2059 956
rect 2348 7457 2859 7630
rect 2348 6709 2378 7457
rect 2834 6709 2859 7457
rect 2348 6506 2859 6709
rect 2858 6449 2859 6506
rect 2348 4878 2859 6449
rect 2858 4821 2859 4878
rect 2348 3250 2859 4821
rect 2858 3193 2859 3250
rect 2348 1622 2859 3193
rect 2858 1565 2859 1622
rect 2348 820 2859 1565
rect 3148 6717 3659 7630
rect 3148 6591 3158 6717
rect 3642 6591 3659 6717
rect 3148 5768 3659 6591
rect 3148 5202 3178 5768
rect 3634 5202 3659 5768
rect 3148 5094 3659 5202
rect 3148 4968 3162 5094
rect 3646 4968 3659 5094
rect 3148 3460 3659 4968
rect 3148 3334 3160 3460
rect 3644 3334 3659 3460
rect 3148 1832 3659 3334
rect 3148 1706 3158 1832
rect 3642 1706 3659 1832
rect 3148 820 3659 1706
rect 4376 7344 4434 7354
rect 4376 346 4434 7111
rect 4496 7024 4554 8171
rect 4496 6780 4554 6791
rect 4616 8094 4674 8095
rect 33764 8094 38644 8242
rect 4616 8018 38644 8094
rect 4496 5495 4554 5517
rect 4496 2460 4554 5262
rect 4616 4106 4674 8018
rect 33764 8010 38644 8018
rect 39091 8010 45075 8242
rect 45169 8010 45603 8242
rect 39091 7970 39156 8010
rect 4736 7905 39156 7970
rect 4736 7344 4794 7905
rect 5108 7753 33185 7847
rect 5108 7701 19892 7753
rect 33067 7701 33185 7753
rect 5108 7609 33185 7701
rect 33426 7609 45886 7847
rect 4982 7498 33435 7512
rect 4982 7294 4999 7498
rect 5136 7294 33435 7498
rect 4982 7278 33435 7294
rect 4736 7098 4794 7111
rect 19586 6278 27923 6512
rect 28159 6278 45886 6512
rect 33202 6277 33433 6278
rect 5747 6215 6173 6226
rect 5747 6067 5761 6215
rect 6157 6067 6173 6215
rect 5747 6055 6173 6067
rect 4932 5883 5150 5902
rect 4932 5880 5019 5883
rect 4932 4243 4956 5880
rect 5128 5172 5150 5883
rect 8078 5495 45886 5508
rect 8078 5487 45221 5495
rect 5128 4785 5443 5172
rect 4932 4240 5019 4243
rect 5128 4240 5150 4785
rect 8078 4501 8099 5487
rect 4932 4219 5150 4240
rect 5278 4367 5389 4371
rect 5278 4360 5651 4367
rect 5002 4218 5149 4219
rect 5278 4138 5285 4360
rect 5381 4356 5651 4360
rect 5381 4141 5566 4356
rect 5639 4141 5651 4356
rect 7843 4292 8099 4501
rect 8287 5288 45221 5487
rect 45595 5288 45886 5495
rect 8287 5274 45886 5288
rect 8287 4292 8312 5274
rect 7843 4269 8312 4292
rect 45101 4236 45404 4320
rect 45770 4236 45886 4320
rect 5381 4138 5651 4141
rect 5278 4131 5651 4138
rect 5278 4127 5389 4131
rect 4616 3849 4674 3873
rect 33053 3824 33063 4062
rect 33115 3824 33186 4062
rect 33427 4043 34526 4062
rect 33427 3959 33565 4043
rect 45101 3959 45404 4043
rect 45770 3959 45886 4043
rect 33427 3824 34526 3959
rect 8196 2800 45886 3038
rect 4496 2402 4674 2460
rect 4496 2229 4554 2249
rect 4496 465 4554 1996
rect 4616 572 4674 2402
rect 4775 2161 5211 2181
rect 4775 641 5042 2161
rect 5198 641 5211 2161
rect 5548 1308 19541 1546
rect 19593 1308 19653 1546
rect 19705 1308 33186 1546
rect 33427 1308 33437 1546
rect 19641 1189 19761 1198
rect 19641 776 19652 1189
rect 19748 776 19761 1189
rect 19641 766 19761 776
rect 32998 1190 33107 1198
rect 32998 776 33009 1190
rect 33096 776 33107 1190
rect 33175 1066 33437 1308
rect 33175 828 45886 1066
rect 32998 766 33107 776
rect 4775 622 5211 641
rect 5426 664 34849 716
rect 5426 572 5478 664
rect 34797 619 34849 664
rect 4616 520 5478 572
rect 5557 563 34367 619
rect 5557 465 5613 563
rect 4496 409 5613 465
rect 33157 431 34367 563
rect 34797 433 45078 619
rect 45486 486 45886 619
rect 34801 431 45078 433
rect 45159 431 45886 486
rect 4376 291 6018 346
rect 5963 116 6018 291
rect 33597 175 33783 363
rect 33983 175 34207 363
rect 34379 175 34391 363
rect 34500 175 44951 363
rect 45159 116 45214 431
rect 45293 350 45599 363
rect 45293 187 45307 350
rect 45581 187 45599 350
rect 45293 175 45599 187
rect 5963 61 45214 116
<< via2 >>
rect 33721 8317 33927 8549
rect 38920 8326 38989 8539
rect 39454 8326 39523 8539
rect 39988 8326 40057 8539
rect 40522 8326 40591 8539
rect 41056 8326 41125 8539
rect 41590 8326 41659 8539
rect 42124 8326 42193 8539
rect 42658 8326 42727 8539
rect 43192 8326 43261 8539
rect 43726 8326 43795 8539
rect 44260 8326 44329 8539
rect 44794 8326 44863 8539
rect 45318 8332 45595 8535
rect 1582 1489 2027 2096
rect 2378 6709 2834 7457
rect 3178 5202 3634 5768
rect 33185 7609 33426 7847
rect 5761 6067 6157 6215
rect 4956 4243 5019 5880
rect 5019 4243 5128 5880
rect 5285 4138 5381 4360
rect 8099 4292 8287 5487
rect 45221 5288 45595 5495
rect 33564 4236 45101 4320
rect 45404 4236 45770 4320
rect 33186 3824 33427 4062
rect 33565 3959 45101 4043
rect 45404 3959 45770 4043
rect 5042 641 5098 2161
rect 33186 1308 33427 1546
rect 19652 776 19748 1189
rect 33009 776 33096 1190
rect 33783 175 33983 363
rect 34391 175 34500 363
rect 45307 187 45581 350
<< metal3 >>
rect 33709 8549 33938 8863
rect 33709 8317 33721 8549
rect 33927 8317 33938 8549
rect 33709 8307 33938 8317
rect 38574 8539 44904 8545
rect 38574 8326 38920 8539
rect 38989 8326 39454 8539
rect 39523 8326 39988 8539
rect 40057 8326 40522 8539
rect 40591 8326 41056 8539
rect 41125 8326 41590 8539
rect 41659 8326 42124 8539
rect 42193 8326 42658 8539
rect 42727 8326 43192 8539
rect 43261 8326 43726 8539
rect 43795 8326 44260 8539
rect 44329 8326 44794 8539
rect 44863 8326 44904 8539
rect 38574 8314 44904 8326
rect 45203 8535 45609 8549
rect 45203 8332 45318 8535
rect 45595 8332 45609 8535
rect 45203 8317 45609 8332
rect 38574 8246 38805 8314
rect 11062 8015 38805 8246
rect 5231 7918 5389 7937
rect 2351 7457 2856 7476
rect 2351 6709 2378 7457
rect 2834 6709 2856 7457
rect 5231 7353 5246 7918
rect 5369 7353 5389 7918
rect 5231 7337 5389 7353
rect 2351 6673 2856 6709
rect 5278 6226 5389 7337
rect 11062 7909 11293 8015
rect 11062 7685 11078 7909
rect 11274 7685 11293 7909
rect 7205 6283 8313 6311
rect 5278 6215 6173 6226
rect 5278 6067 5761 6215
rect 6157 6067 6173 6215
rect 7205 6100 7254 6283
rect 7704 6100 8313 6283
rect 7205 6074 8313 6100
rect 5278 6055 6173 6067
rect 4932 5880 5150 5902
rect 3150 5768 3654 5800
rect 3150 5202 3178 5768
rect 3634 5202 3654 5768
rect 3150 5176 3654 5202
rect 4932 4243 4956 5880
rect 5128 4243 5150 5880
rect 4932 4219 5150 4243
rect 5278 4360 5389 6055
rect 8076 5487 8313 6074
rect 5278 4138 5285 4360
rect 5381 4138 5389 4360
rect 4675 2161 5111 2181
rect 1552 2096 2057 2126
rect 1552 1489 1582 2096
rect 2027 1489 2057 2096
rect 1552 1461 2057 1489
rect 4675 641 4942 2161
rect 5098 641 5111 2161
rect 5278 981 5389 4138
rect 8076 4292 8099 5487
rect 8287 4292 8313 5487
rect 8076 2233 8313 4292
rect 7221 2202 8313 2233
rect 7221 2019 7266 2202
rect 7716 2019 8313 2202
rect 7221 1996 8313 2019
rect 4675 622 5111 641
rect 5232 960 5390 981
rect 5232 395 5246 960
rect 5369 395 5390 960
rect 5232 381 5390 395
rect 11062 634 11293 7685
rect 33175 7847 33437 7855
rect 33175 7609 33185 7847
rect 33426 7609 33437 7847
rect 33175 4062 33437 7609
rect 45203 5508 45322 8317
rect 45203 5495 45615 5508
rect 45203 5288 45221 5495
rect 45595 5288 45615 5495
rect 45203 5274 45615 5288
rect 33539 4409 45113 4454
rect 33539 4236 33564 4409
rect 45101 4236 45113 4409
rect 33539 4220 45113 4236
rect 33175 3824 33186 4062
rect 33427 4043 45113 4062
rect 33427 3870 33521 4043
rect 45101 3870 45113 4043
rect 33427 3824 45113 3870
rect 33175 1546 33437 3824
rect 33175 1308 33186 1546
rect 33427 1308 33437 1546
rect 33175 1295 33437 1308
rect 11062 397 11079 634
rect 11277 397 11293 634
rect 11062 383 11293 397
rect 19641 1189 19761 1198
rect 19641 776 19652 1189
rect 19748 776 19761 1189
rect 19641 25 19761 776
rect 32998 1190 33107 1198
rect 32998 776 33009 1190
rect 33096 776 33107 1190
rect 32998 607 33107 776
rect 32998 498 34500 607
rect 33776 363 33991 385
rect 34391 369 34500 498
rect 33776 175 33783 363
rect 33983 175 33991 363
rect 33776 0 33991 175
rect 34384 363 34506 369
rect 34384 175 34391 363
rect 34500 175 34506 363
rect 34384 169 34506 175
rect 45203 363 45322 5274
rect 45392 4409 45903 4454
rect 45392 4236 45404 4409
rect 45770 4236 45903 4409
rect 45392 4220 45903 4236
rect 45392 4043 45903 4062
rect 45392 3870 45404 4043
rect 45770 3870 45903 4043
rect 45392 3824 45903 3870
rect 45203 350 45599 363
rect 45203 187 45307 350
rect 45581 187 45599 350
rect 45203 174 45599 187
<< via3 >>
rect 2378 6709 2834 7457
rect 5246 7353 5369 7918
rect 11078 7685 11274 7909
rect 7254 6100 7704 6283
rect 3178 5202 3634 5768
rect 4956 4243 5128 5880
rect 7112 4802 7851 5156
rect 1582 1489 2027 2096
rect 4942 641 5042 2161
rect 5042 641 5098 2161
rect 7204 3165 7930 3501
rect 7266 2019 7716 2202
rect 5246 395 5369 960
rect 33564 4320 45101 4409
rect 33564 4236 45101 4320
rect 33521 3959 33565 4043
rect 33565 3959 45101 4043
rect 33521 3870 45101 3959
rect 11079 397 11277 634
rect 45404 4320 45770 4409
rect 45404 4236 45770 4320
rect 45404 3959 45770 4043
rect 45404 3870 45770 3959
<< metal4 >>
rect 5231 7924 5389 7937
rect 5231 7918 5625 7924
rect 1098 7457 4102 7504
rect 1098 6709 2378 7457
rect 2834 6709 4102 7457
rect 5231 7353 5246 7918
rect 5369 7820 5625 7918
rect 10789 7909 11293 7924
rect 10789 7821 11078 7909
rect 5369 7353 5389 7820
rect 11062 7685 11078 7821
rect 11274 7685 11293 7909
rect 11062 7668 11293 7685
rect 5231 7337 5389 7353
rect 1098 6104 4102 6709
rect 7410 6311 7540 6688
rect 7223 6283 7739 6311
rect 7223 6100 7254 6283
rect 7704 6100 7739 6283
rect 7223 6074 7739 6100
rect 1098 5880 45903 5902
rect 1098 5768 4956 5880
rect 1098 5202 3178 5768
rect 3634 5202 4956 5768
rect 1098 4243 4956 5202
rect 5128 5156 45903 5880
rect 5128 4802 7112 5156
rect 7851 4802 45903 5156
rect 5128 4409 45903 4802
rect 5128 4243 33564 4409
rect 1098 4236 33564 4243
rect 45101 4236 45404 4409
rect 45770 4236 45903 4409
rect 1098 4217 45903 4236
rect 1098 4043 45903 4066
rect 1098 3870 33521 4043
rect 45101 3870 45404 4043
rect 45770 3870 45903 4043
rect 1098 3501 45903 3870
rect 1098 3165 7204 3501
rect 7930 3165 45903 3501
rect 1098 2381 45903 3165
rect 7234 2202 7750 2233
rect 1098 2161 5111 2182
rect 1098 2096 4942 2161
rect 1098 1489 1582 2096
rect 2027 1489 4942 2096
rect 1098 641 4942 1489
rect 5098 641 5111 2161
rect 7234 2019 7266 2202
rect 7716 2019 7750 2202
rect 7234 1996 7750 2019
rect 7423 1620 7553 1996
rect 1098 622 5111 641
rect 5232 960 5390 981
rect 5232 395 5246 960
rect 5369 487 5390 960
rect 11062 634 11293 649
rect 11062 487 11079 634
rect 5369 395 5634 487
rect 5232 383 5634 395
rect 10810 397 11079 487
rect 11277 397 11293 634
rect 10810 383 11293 397
rect 5232 381 5390 383
use bias_amp  bias_amp_0
timestamp 1717075507
transform 1 0 0 0 1 0
box 5361 2480 8196 5306
use bias_nstack  bias_nstack_0
array 0 22 -534 0 0 -3895
timestamp 1717035242
transform -1 0 37396 0 -1 1202
box 3258 -2860 3926 1035
use bias_pstack  bias_pstack_0
array 0 22 534 0 0 -4355
timestamp 1717035242
transform 1 0 31443 0 -1 4608
box 1986 -3967 2714 388
use sky130_fd_pr__cap_mim_m3_1_MQZGVK  sky130_fd_pr__cap_mim_m3_1_MQZGVK_0 paramcells
timestamp 1717035242
transform 0 1 8149 1 0 7238
box -686 -2640 686 2640
use sky130_fd_pr__cap_mim_m3_1_MQZGVK  sky130_fd_pr__cap_mim_m3_1_MQZGVK_1
timestamp 1717035242
transform 0 1 8170 -1 0 1069
box -686 -2640 686 2640
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  sky130_fd_pr__diode_pw2nd_05v5_FT76RJ_0 paramcells
timestamp 1717075507
transform 1 0 6054 0 1 5446
box -183 -183 183 183
use sky130_fd_pr__res_high_po_0p35_L4QTBM  sky130_fd_pr__res_high_po_0p35_L4QTBM_0 paramcells
timestamp 1717035242
transform 1 0 13944 0 1 4182
box -5679 -3582 5679 3582
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform 1 0 3486 0 1 4217
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_1
timestamp 1715205430
transform 1 0 3486 0 1 961
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_2
timestamp 1715205430
transform 1 0 3486 0 1 2589
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_3
timestamp 1715205430
transform 1 0 3486 0 -1 5845
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_4
timestamp 1715205430
transform 1 0 3486 0 1 5845
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_11
timestamp 1715205430
transform 1 0 3486 0 -1 2589
box -66 -43 450 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform 1 0 3870 0 1 4217
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_1
timestamp 1715205430
transform 1 0 3870 0 -1 2589
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_2
timestamp 1715205430
transform 1 0 3870 0 1 2589
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_3
timestamp 1715205430
transform 1 0 3870 0 -1 5845
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_4
timestamp 1715205430
transform 1 0 3870 0 1 5845
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_11
timestamp 1715205430
transform 1 0 3870 0 1 961
box -66 -43 162 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_2 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform 1 0 3486 0 -1 4217
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_4
timestamp 1715205430
transform 1 0 3486 0 -1 7473
box -66 -43 546 897
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
array 0 0 2592 0 3 1628
timestamp 1715205430
transform 1 0 1374 0 1 961
box -66 -43 2178 1671
use sky130_fd_pr__res_high_po_0p35_P35QVK  XR2 paramcells
timestamp 1717035242
transform 1 0 26381 0 1 4182
box -6758 -3582 6758 3582
<< labels >>
flabel metal3 33776 0 33991 153 0 FreeSans 1600 90 0 0 snk_test0
port 40 nsew
flabel metal3 33709 8630 33938 8863 0 FreeSans 1600 90 0 0 src_test0
port 45 nsew
flabel metal1 1072 6185 1472 6253 0 FreeSans 480 0 0 0 ref_sel_vbg
port 52 nsew
flabel metal1 1072 4557 1472 4625 0 FreeSans 480 0 0 0 ena
port 53 nsew
flabel metal1 1072 2929 1472 2997 0 FreeSans 480 0 0 0 ena_src_test0
port 61 nsew
flabel metal1 1072 1301 1472 1369 0 FreeSans 480 0 0 0 ena_snk_test0
port 60 nsew
flabel metal1 4150 3892 4150 3892 0 FreeSans 480 0 0 0 enb_test0_3v3
flabel metal1 4127 5281 4127 5281 0 FreeSans 480 0 0 0 ena_3v3
flabel metal1 4118 6906 4118 6906 0 FreeSans 480 0 0 0 ena_vbg_3v3
flabel metal1 4133 7133 4133 7133 0 FreeSans 480 0 0 0 enb_vbg_3v3
flabel metal1 5441 8326 5562 8557 0 FreeSans 1600 90 0 0 vbg
port 56 nsew
flabel metal2 32539 7935 32539 7935 0 FreeSans 640 0 0 0 enb_vbg_3v3
flabel metal2 32553 8052 32553 8052 0 FreeSans 640 0 0 0 enb_test0_3v3
flabel metal2 32634 592 32634 592 0 FreeSans 640 0 0 0 ena_test0_3v3
flabel space 32658 693 32658 693 0 FreeSans 640 0 0 0 ena_3v3
flabel metal3 19641 25 19761 381 0 FreeSans 1600 90 0 0 ref_in
port 57 nsew
flabel metal2 32668 85 32668 85 0 FreeSans 640 0 0 0 enb_vbg_3v3
flabel metal2 32589 8212 32589 8212 0 FreeSans 640 0 0 0 ena_vbg_3v3
flabel metal4 1098 4217 1698 5902 0 FreeSans 3200 90 0 0 avdd
port 59 nsew
flabel metal4 1098 2381 1698 4066 0 FreeSans 3200 90 0 0 avss
port 12 nsew
flabel metal4 1098 6104 1698 7504 0 FreeSans 3200 90 0 0 dvdd
port 58 n
flabel metal4 1098 622 1698 2182 0 FreeSans 3200 90 0 0 dvss
port 50 nsew
flabel metal1 4492 2022 4492 2022 0 FreeSans 480 0 0 0 ena_test0_3v3
<< end >>
