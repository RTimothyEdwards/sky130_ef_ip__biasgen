magic
tech sky130A
magscale 1 2
timestamp 1719420833
<< error_s >>
rect 135078 -10275 135978 -9375
<< dnwell >>
rect 96152 19519 138230 27371
rect 89743 9519 138229 17371
rect 89743 -481 138229 7371
rect 135078 -10481 138229 -2629
<< nwell >>
rect 96043 27165 138339 27480
rect 96043 19725 96358 27165
rect 138024 19725 138339 27165
rect 96043 19410 138339 19725
rect 89634 17165 138338 17480
rect 89634 9725 89949 17165
rect 138023 9725 138338 17165
rect 89634 9410 138338 9725
rect 89634 7165 138338 7480
rect 89634 -275 89949 7165
rect 138023 -275 138338 7165
rect 89634 -590 138338 -275
rect 135078 -2835 138338 -2520
rect 138023 -10275 138338 -2835
rect 135078 -10590 138338 -10275
<< pwell >>
rect 125398 19725 125486 19747
rect 108895 9725 108983 9747
rect 108895 -275 108983 -253
<< mvpsubdiff >>
rect 95923 27570 95983 27604
rect 137413 27570 137603 27604
rect 138399 27570 138459 27604
rect 95923 27544 95957 27570
rect 88137 26982 88197 27016
rect 95249 26982 95309 27016
rect 88137 26956 88171 26982
rect 88137 20052 88171 20078
rect 95275 26956 95309 26982
rect 95275 20052 95309 20078
rect 88137 20018 88197 20052
rect 95249 20018 95309 20052
rect 138425 27544 138459 27570
rect 95923 19298 95957 19324
rect 138425 19298 138459 19324
rect 95923 19264 95983 19298
rect 137413 19264 137603 19298
rect 138399 19264 138459 19298
rect 89514 17570 89574 17604
rect 90370 17570 90560 17604
rect 138398 17570 138458 17604
rect 89514 17544 89548 17570
rect 138424 17544 138458 17570
rect 89514 9298 89548 9324
rect 138424 9298 138458 9324
rect 89514 9264 89574 9298
rect 90370 9264 90560 9298
rect 138398 9264 138458 9298
rect 89514 7570 89574 7604
rect 90370 7570 90560 7604
rect 138398 7570 138458 7604
rect 89514 7544 89548 7570
rect 138424 7544 138458 7570
rect 89514 -702 89548 -676
rect 138424 -702 138458 -676
rect 89514 -736 89574 -702
rect 90370 -736 90560 -702
rect 138398 -736 138458 -702
rect 135144 -2430 135416 -2396
rect 138398 -2430 138458 -2396
rect 138424 -2456 138458 -2430
rect 138424 -10702 138458 -10676
rect 135144 -10736 135416 -10702
rect 138398 -10736 138458 -10702
<< mvnsubdiff >>
rect 96109 27394 138273 27414
rect 96109 27360 96189 27394
rect 137413 27360 137603 27394
rect 138193 27360 138273 27394
rect 96109 27340 138273 27360
rect 96109 27334 96183 27340
rect 96109 19556 96129 27334
rect 96163 19556 96183 27334
rect 96109 19550 96183 19556
rect 138199 27334 138273 27340
rect 138199 19556 138219 27334
rect 138253 19556 138273 27334
rect 138199 19550 138273 19556
rect 96109 19530 138273 19550
rect 96109 19496 96189 19530
rect 137413 19496 137603 19530
rect 138193 19496 138273 19530
rect 96109 19476 138273 19496
rect 89700 17394 138272 17414
rect 89700 17360 89780 17394
rect 90370 17360 90560 17394
rect 138192 17360 138272 17394
rect 89700 17340 138272 17360
rect 89700 17334 89774 17340
rect 89700 9556 89720 17334
rect 89754 9556 89774 17334
rect 89700 9550 89774 9556
rect 138198 17334 138272 17340
rect 138198 9556 138218 17334
rect 138252 9556 138272 17334
rect 138198 9550 138272 9556
rect 89700 9530 138272 9550
rect 89700 9496 89780 9530
rect 90370 9496 90560 9530
rect 138192 9496 138272 9530
rect 89700 9476 138272 9496
rect 89700 7394 138272 7414
rect 89700 7360 89780 7394
rect 90370 7360 90560 7394
rect 138192 7360 138272 7394
rect 89700 7340 138272 7360
rect 89700 7334 89774 7340
rect 89700 -444 89720 7334
rect 89754 -444 89774 7334
rect 89700 -450 89774 -444
rect 138198 7334 138272 7340
rect 138198 -444 138218 7334
rect 138252 -444 138272 7334
rect 138198 -450 138272 -444
rect 89700 -470 138272 -450
rect 89700 -504 89780 -470
rect 90370 -504 90560 -470
rect 138192 -504 138272 -470
rect 89700 -524 138272 -504
rect 135144 -2606 138272 -2586
rect 135144 -2640 135416 -2606
rect 138192 -2640 138272 -2606
rect 135144 -2660 138272 -2640
rect 138198 -2666 138272 -2660
rect 138198 -10444 138218 -2666
rect 138252 -10444 138272 -2666
rect 138198 -10450 138272 -10444
rect 135144 -10470 138272 -10450
rect 135144 -10504 135416 -10470
rect 138192 -10504 138272 -10470
rect 135144 -10524 138272 -10504
<< mvpsubdiffcont >>
rect 95983 27570 137413 27604
rect 137603 27570 138399 27604
rect 88197 26982 95249 27016
rect 88137 20078 88171 26956
rect 95275 20078 95309 26956
rect 88197 20018 95249 20052
rect 95923 19324 95957 27544
rect 138425 19324 138459 27544
rect 95983 19264 137413 19298
rect 137603 19264 138399 19298
rect 89574 17570 90370 17604
rect 90560 17570 138398 17604
rect 89514 9324 89548 17544
rect 138424 9324 138458 17544
rect 89574 9264 90370 9298
rect 90560 9264 138398 9298
rect 89574 7570 90370 7604
rect 90560 7570 138398 7604
rect 89514 -676 89548 7544
rect 138424 -676 138458 7544
rect 89574 -736 90370 -702
rect 90560 -736 138398 -702
rect 135416 -2430 138398 -2396
rect 138424 -10676 138458 -2456
rect 135416 -10736 138398 -10702
<< mvnsubdiffcont >>
rect 96189 27360 137413 27394
rect 137603 27360 138193 27394
rect 96129 19556 96163 27334
rect 138219 19556 138253 27334
rect 96189 19496 137413 19530
rect 137603 19496 138193 19530
rect 89780 17360 90370 17394
rect 90560 17360 138192 17394
rect 89720 9556 89754 17334
rect 138218 9556 138252 17334
rect 89780 9496 90370 9530
rect 90560 9496 138192 9530
rect 89780 7360 90370 7394
rect 90560 7360 138192 7394
rect 89720 -444 89754 7334
rect 138218 -444 138252 7334
rect 89780 -504 90370 -470
rect 90560 -504 138192 -470
rect 135416 -2640 138192 -2606
rect 138218 -10444 138252 -2666
rect 135416 -10504 138192 -10470
<< locali >>
rect 95923 27570 95983 27604
rect 137413 27570 137603 27604
rect 138399 27570 138459 27604
rect 95923 27555 138459 27570
rect 95923 27544 95969 27555
rect 88137 26982 88197 27016
rect 95249 26982 95923 27016
rect 88137 26956 95923 26982
rect 88171 26894 95275 26956
rect 88171 20140 88265 26894
rect 91871 26394 91918 26460
rect 90110 25566 90280 25582
rect 90110 25464 90131 25566
rect 90264 25464 90280 25566
rect 90110 25448 90280 25464
rect 92702 25566 92872 25582
rect 92702 25464 92723 25566
rect 92856 25464 92872 25566
rect 92702 25448 92872 25464
rect 91871 24766 91918 24832
rect 90110 23938 90280 23954
rect 90110 23836 90131 23938
rect 90264 23836 90280 23938
rect 90110 23820 90280 23836
rect 92702 23938 92872 23954
rect 92702 23836 92723 23938
rect 92856 23836 92872 23938
rect 92702 23820 92872 23836
rect 91871 23138 91918 23204
rect 90110 22310 90280 22326
rect 90110 22208 90131 22310
rect 90264 22208 90280 22310
rect 90110 22192 90280 22208
rect 92702 22310 92872 22326
rect 92702 22208 92723 22310
rect 92856 22208 92872 22310
rect 92702 22192 92872 22208
rect 91871 21510 91918 21576
rect 90110 20682 90280 20698
rect 90110 20580 90131 20682
rect 90264 20580 90280 20682
rect 90110 20564 90280 20580
rect 92702 20682 92872 20698
rect 92702 20580 92723 20682
rect 92856 20580 92872 20682
rect 92702 20564 92872 20580
rect 95192 20140 95275 26894
rect 88171 20078 95275 20140
rect 95309 26819 95923 26956
rect 95309 20078 95923 20214
rect 88137 20052 95923 20078
rect 88137 20018 88197 20052
rect 95249 20018 95923 20052
rect 95220 20017 95923 20018
rect 95957 19324 95969 27544
rect 95923 19314 95969 19324
rect 96021 27471 138361 27555
rect 96021 19410 96065 27471
rect 96129 27360 96189 27394
rect 137413 27360 137603 27394
rect 138193 27360 138253 27394
rect 96129 27334 138253 27360
rect 96163 27329 138219 27334
rect 96163 19556 96194 27329
rect 96129 19552 96194 19556
rect 96253 27292 138129 27329
rect 96253 27226 96850 27292
rect 97000 27226 138129 27292
rect 96253 27175 138129 27226
rect 96253 19709 96300 27175
rect 138082 19709 138129 27175
rect 96253 19552 138129 19709
rect 138188 19556 138219 27329
rect 138188 19552 138253 19556
rect 96129 19530 138253 19552
rect 96129 19496 96189 19530
rect 137413 19496 137603 19530
rect 138193 19496 138253 19530
rect 138317 19410 138361 27471
rect 96021 19323 138361 19410
rect 96021 19314 96074 19323
rect 95923 19298 96074 19314
rect 95923 19264 95983 19298
rect 137413 19264 137603 19323
rect 138308 19314 138361 19323
rect 138413 27544 138459 27555
rect 138413 19324 138425 27544
rect 138459 26819 138541 27016
rect 138459 20017 138541 20214
rect 138413 19314 138459 19324
rect 138308 19298 138459 19314
rect 138399 19264 138459 19298
rect 89514 17570 89574 17604
rect 90370 17570 90560 17604
rect 138398 17570 138458 17604
rect 89514 17555 138458 17570
rect 89514 17544 89560 17555
rect 89432 16819 89514 17016
rect 89432 10017 89514 10214
rect 89548 9324 89560 17544
rect 89514 9314 89560 9324
rect 89612 17471 138360 17555
rect 89612 9410 89656 17471
rect 89720 17360 89780 17394
rect 90370 17360 90560 17394
rect 138192 17360 138252 17394
rect 89720 17334 138252 17360
rect 89754 17329 138218 17334
rect 89754 9556 89785 17329
rect 89720 9552 89785 9556
rect 89844 17292 138128 17329
rect 89844 17226 137381 17292
rect 137531 17226 138128 17292
rect 89844 17175 138128 17226
rect 89844 9709 89891 17175
rect 138081 9709 138128 17175
rect 89844 9552 138128 9709
rect 138187 9556 138218 17329
rect 138187 9552 138252 9556
rect 89720 9530 138252 9552
rect 89720 9496 89780 9530
rect 90370 9496 90560 9530
rect 138192 9496 138252 9530
rect 138316 9410 138360 17471
rect 89612 9323 138360 9410
rect 89612 9314 89665 9323
rect 89514 9298 89665 9314
rect 89514 9264 89574 9298
rect 90370 9264 90560 9323
rect 138307 9314 138360 9323
rect 138412 17544 138458 17555
rect 138412 9324 138424 17544
rect 138458 16819 138540 17016
rect 138458 10017 138540 10214
rect 138412 9314 138458 9324
rect 138307 9298 138458 9314
rect 138398 9264 138458 9298
rect 89514 7570 89574 7604
rect 90370 7570 90560 7604
rect 138398 7570 138458 7604
rect 89514 7555 138458 7570
rect 89514 7544 89560 7555
rect 89432 6819 89514 7016
rect 89432 17 89514 214
rect 89548 -676 89560 7544
rect 89514 -686 89560 -676
rect 89612 7471 138360 7555
rect 89612 -590 89656 7471
rect 89720 7360 89780 7394
rect 90370 7360 90560 7394
rect 138192 7360 138252 7394
rect 89720 7334 138252 7360
rect 89754 7329 138218 7334
rect 89754 -444 89785 7329
rect 89720 -448 89785 -444
rect 89844 7292 138128 7329
rect 89844 7226 137381 7292
rect 137531 7226 138128 7292
rect 89844 7175 138128 7226
rect 89844 -291 89891 7175
rect 138081 -291 138128 7175
rect 89844 -448 138128 -291
rect 138187 -444 138218 7329
rect 138187 -448 138252 -444
rect 89720 -470 138252 -448
rect 89720 -504 89780 -470
rect 90370 -504 90560 -470
rect 138192 -504 138252 -470
rect 138316 -590 138360 7471
rect 89612 -677 138360 -590
rect 89612 -686 89665 -677
rect 89514 -702 89665 -686
rect 89514 -736 89574 -702
rect 90370 -736 90560 -677
rect 138307 -686 138360 -677
rect 138412 7544 138458 7555
rect 138412 -676 138424 7544
rect 138458 6819 138540 7016
rect 138458 17 138540 214
rect 138412 -686 138458 -676
rect 138307 -702 138458 -686
rect 138398 -736 138458 -702
rect 135144 -2430 135416 -2396
rect 138398 -2430 138458 -2396
rect 135144 -2445 138458 -2430
rect 135144 -2529 138360 -2445
rect 135152 -2640 135416 -2606
rect 138192 -2640 138252 -2606
rect 135152 -2666 138252 -2640
rect 135152 -2671 138218 -2666
rect 135152 -2825 138128 -2671
rect 138081 -10291 138128 -2825
rect 135144 -10448 138128 -10291
rect 138187 -10444 138218 -2671
rect 138187 -10448 138252 -10444
rect 135144 -10470 138252 -10448
rect 135144 -10504 135416 -10470
rect 138192 -10504 138252 -10470
rect 138316 -10590 138360 -2529
rect 135144 -10677 138360 -10590
rect 135144 -10736 135416 -10677
rect 138307 -10686 138360 -10677
rect 138412 -2456 138458 -2445
rect 138412 -10676 138424 -2456
rect 138458 -3181 138540 -2984
rect 138458 -9983 138540 -9786
rect 138412 -10686 138458 -10676
rect 138307 -10702 138458 -10686
rect 138398 -10736 138458 -10702
<< viali >>
rect 89614 26424 89660 26603
rect 92206 26424 92252 26603
rect 94415 26116 94463 26347
rect 90131 25464 90264 25566
rect 92723 25464 92856 25566
rect 89614 24796 89660 24975
rect 92206 24796 92252 24975
rect 94415 24488 94463 24719
rect 90131 23836 90264 23938
rect 92723 23836 92856 23938
rect 89614 23168 89660 23347
rect 92206 23168 92252 23347
rect 94415 22860 94463 23091
rect 90131 22208 90264 22310
rect 92723 22208 92856 22310
rect 89614 21540 89660 21719
rect 92206 21540 92252 21719
rect 94415 21232 94463 21463
rect 90131 20580 90264 20682
rect 92723 20580 92856 20682
rect 95969 19314 96021 27555
rect 96194 19552 96253 27329
rect 96850 27226 97000 27292
rect 138129 19552 138188 27329
rect 96074 19298 137413 19323
rect 96074 19279 137413 19298
rect 137603 19298 138308 19323
rect 138361 19314 138413 27555
rect 137603 19279 138308 19298
rect 89560 9314 89612 17555
rect 89785 9552 89844 17329
rect 137381 17226 137531 17292
rect 138128 9552 138187 17329
rect 89665 9298 90370 9323
rect 89665 9279 90370 9298
rect 90560 9298 138307 9323
rect 138360 9314 138412 17555
rect 90560 9279 138307 9298
rect 89560 -686 89612 7555
rect 89785 -448 89844 7329
rect 137381 7226 137531 7292
rect 138128 -448 138187 7329
rect 89665 -702 90370 -677
rect 89665 -721 90370 -702
rect 90560 -702 138307 -677
rect 138360 -686 138412 7555
rect 90560 -721 138307 -702
rect 138128 -10448 138187 -2671
rect 135416 -10702 138307 -10677
rect 138360 -10686 138412 -2445
rect 135416 -10721 138307 -10702
<< metal1 >>
rect 95933 27555 96049 27597
rect 88353 26831 95047 26845
rect 88353 26672 93083 26831
rect 94358 26672 95047 26831
rect 89605 26614 89669 26616
rect 92201 26615 92265 26616
rect 89605 26414 89611 26614
rect 89663 26414 89669 26614
rect 89605 26412 89669 26414
rect 92200 26614 92265 26615
rect 92200 26603 92207 26614
rect 92200 26424 92206 26603
rect 92200 26414 92207 26424
rect 92259 26414 92265 26614
rect 92200 26412 92259 26414
rect 89613 26400 89653 26412
rect 92201 26329 92241 26412
rect 94414 26384 95669 26424
rect 94414 26353 94454 26384
rect 94399 26347 94475 26353
rect 94399 26116 94415 26347
rect 94463 26116 94475 26347
rect 95663 26224 95669 26384
rect 95721 26224 95727 26424
rect 94399 26110 94475 26116
rect 88364 25866 90501 26039
rect 91780 25866 95047 26039
rect 88811 25746 88829 25803
rect 89205 25746 95047 25803
rect 90110 25566 90280 25582
rect 90110 25464 90131 25566
rect 90264 25464 90280 25566
rect 90110 25448 90280 25464
rect 92702 25566 92872 25582
rect 92702 25464 92723 25566
rect 92856 25464 92872 25566
rect 92702 25448 92872 25464
rect 88364 25049 93085 25222
rect 94355 25049 95047 25222
rect 89608 24986 89667 24987
rect 92199 24986 92265 24988
rect 89605 24786 89611 24986
rect 89663 24786 89669 24986
rect 92199 24975 92207 24986
rect 92199 24796 92206 24975
rect 92199 24786 92207 24796
rect 92259 24786 92265 24986
rect 89605 24784 89669 24786
rect 92200 24784 92259 24786
rect 89613 24780 89653 24784
rect 92201 24701 92241 24784
rect 94414 24756 95563 24796
rect 94414 24725 94454 24756
rect 94399 24719 94475 24725
rect 94399 24488 94415 24719
rect 94463 24488 94475 24719
rect 95557 24596 95563 24756
rect 95615 24596 95621 24796
rect 94399 24482 94475 24488
rect 88347 24238 90505 24411
rect 91784 24238 95047 24411
rect 88811 24118 88825 24175
rect 89205 24118 95047 24175
rect 90110 23938 90280 23954
rect 90110 23836 90131 23938
rect 90264 23836 90280 23938
rect 90110 23820 90280 23836
rect 92702 23938 92872 23954
rect 92702 23836 92723 23938
rect 92856 23836 92872 23938
rect 92702 23820 92872 23836
rect 88375 23422 93087 23595
rect 94357 23422 95047 23595
rect 92201 23359 92265 23360
rect 89608 23358 89667 23359
rect 92200 23358 92265 23359
rect 89605 23158 89611 23358
rect 89663 23158 89669 23358
rect 89605 23156 89669 23158
rect 92200 23347 92207 23358
rect 92200 23168 92206 23347
rect 92259 23328 92265 23358
rect 92200 23158 92207 23168
rect 92259 23158 92265 23288
rect 92200 23156 92259 23158
rect 89613 23150 89653 23156
rect 94414 23128 95481 23168
rect 94414 23097 94454 23128
rect 94399 23091 94475 23097
rect 94399 22860 94415 23091
rect 94463 22860 94475 23091
rect 95475 22968 95481 23128
rect 95533 22968 95539 23168
rect 94399 22854 94475 22860
rect 88358 22622 90501 22795
rect 91780 22622 95047 22795
rect 88811 22490 88822 22547
rect 89205 22490 95047 22547
rect 90110 22310 90280 22326
rect 90110 22208 90131 22310
rect 90264 22208 90280 22310
rect 90110 22192 90280 22208
rect 92702 22310 92872 22326
rect 92702 22208 92723 22310
rect 92856 22208 92872 22310
rect 92702 22192 92872 22208
rect 88391 21800 93083 21973
rect 94353 21800 95047 21973
rect 89608 21730 89667 21731
rect 92199 21730 92265 21732
rect 89605 21530 89611 21730
rect 89663 21530 89669 21730
rect 92199 21719 92207 21730
rect 92199 21540 92206 21719
rect 92259 21700 92265 21730
rect 92199 21530 92207 21540
rect 92259 21530 92265 21660
rect 89605 21528 89669 21530
rect 92200 21528 92259 21530
rect 89613 21510 89653 21528
rect 94418 21500 95391 21540
rect 94418 21469 94458 21500
rect 94402 21463 94475 21469
rect 94402 21232 94415 21463
rect 94463 21232 94475 21463
rect 95385 21340 95391 21500
rect 95443 21340 95449 21540
rect 95933 21312 95969 27555
rect 94402 21226 94475 21232
rect 95759 21281 95969 21312
rect 88347 20983 90501 21156
rect 91780 20983 95047 21156
rect 88811 20862 88822 20919
rect 89205 20862 95047 20919
rect 90110 20682 90280 20698
rect 90110 20580 90131 20682
rect 90264 20580 90280 20682
rect 90110 20564 90280 20580
rect 92702 20682 92872 20698
rect 92702 20580 92723 20682
rect 92856 20580 92872 20682
rect 92702 20564 92872 20580
rect 88425 20261 93088 20339
rect 94360 20261 95047 20339
rect 95759 20142 95788 21281
rect 95759 20110 95969 20142
rect 95933 19314 95969 20110
rect 96021 19342 96049 27555
rect 138333 27555 138449 27597
rect 96150 27329 96288 27380
rect 96150 25099 96194 27329
rect 96253 25099 96288 27329
rect 138094 27329 138232 27380
rect 96837 27292 97016 27304
rect 96837 27226 96850 27292
rect 97000 27281 97016 27292
rect 97000 27229 97151 27281
rect 97000 27226 97016 27229
rect 96837 27216 97016 27226
rect 96150 23457 96166 25099
rect 96273 23457 96288 25099
rect 96150 19552 96194 23457
rect 96253 19552 96288 23457
rect 138094 25099 138129 27329
rect 138188 25099 138232 27329
rect 138094 23457 138109 25099
rect 138216 23457 138232 25099
rect 96150 19505 96288 19552
rect 97096 19342 97150 19646
rect 138094 19552 138129 23457
rect 138188 19552 138232 23457
rect 138094 19505 138232 19552
rect 138333 19342 138361 27555
rect 138413 21312 138449 27555
rect 138413 21281 138541 21312
rect 96021 19323 138361 19342
rect 96021 19314 96074 19323
rect 95933 19279 96074 19314
rect 137413 19279 137603 19323
rect 138308 19314 138361 19323
rect 138413 20110 138541 20142
rect 138413 19314 138449 20110
rect 138308 19279 138449 19314
rect 95933 19264 138449 19279
rect 89524 17555 89640 17597
rect 89524 11312 89560 17555
rect 89432 11281 89560 11312
rect 89432 10110 89560 10142
rect 89524 9314 89560 10110
rect 89612 9342 89640 17555
rect 138332 17555 138448 17597
rect 89741 17329 89879 17380
rect 89741 15099 89785 17329
rect 89844 15099 89879 17329
rect 138093 17329 138231 17380
rect 137365 17292 137544 17304
rect 137365 17281 137381 17292
rect 137230 17229 137381 17281
rect 137365 17226 137381 17229
rect 137531 17226 137544 17292
rect 137365 17216 137544 17226
rect 89741 13457 89757 15099
rect 89864 13457 89879 15099
rect 89741 9552 89785 13457
rect 89844 9552 89879 13457
rect 138093 15099 138128 17329
rect 138187 15099 138231 17329
rect 138093 13457 138108 15099
rect 138215 13457 138231 15099
rect 89741 9505 89879 9552
rect 137231 9342 137285 9646
rect 138093 9552 138128 13457
rect 138187 9552 138231 13457
rect 138093 9505 138231 9552
rect 138332 9342 138360 17555
rect 138412 11312 138448 17555
rect 138412 11281 138540 11312
rect 89612 9323 138360 9342
rect 89612 9314 89665 9323
rect 89524 9279 89665 9314
rect 90370 9279 90560 9323
rect 138307 9314 138360 9323
rect 138412 10110 138540 10142
rect 138412 9314 138448 10110
rect 138307 9279 138448 9314
rect 89524 9264 138448 9279
rect 89524 7555 89640 7597
rect 89524 1312 89560 7555
rect 89432 1281 89560 1312
rect 89432 110 89560 142
rect 89524 -686 89560 110
rect 89612 -658 89640 7555
rect 138332 7555 138448 7597
rect 89741 7329 89879 7380
rect 89741 5099 89785 7329
rect 89844 5099 89879 7329
rect 138093 7329 138231 7380
rect 137365 7292 137544 7304
rect 137365 7281 137381 7292
rect 137230 7229 137381 7281
rect 137365 7226 137381 7229
rect 137531 7226 137544 7292
rect 137365 7216 137544 7226
rect 89741 3457 89757 5099
rect 89864 3457 89879 5099
rect 89741 -448 89785 3457
rect 89844 -448 89879 3457
rect 138093 5099 138128 7329
rect 138187 5099 138231 7329
rect 138093 3457 138108 5099
rect 138215 3457 138231 5099
rect 89741 -495 89879 -448
rect 137231 -658 137285 -354
rect 138093 -448 138128 3457
rect 138187 -448 138231 3457
rect 138093 -495 138231 -448
rect 138332 -658 138360 7555
rect 138412 1312 138448 7555
rect 138412 1281 138540 1312
rect 89612 -677 138360 -658
rect 89612 -686 89665 -677
rect 89524 -721 89665 -686
rect 90370 -721 90560 -677
rect 138307 -686 138360 -677
rect 138412 110 138540 142
rect 138412 -686 138448 110
rect 138307 -721 138448 -686
rect 89524 -736 138448 -721
rect 138332 -2445 138448 -2403
rect 138093 -2671 138231 -2620
rect 138093 -4901 138128 -2671
rect 138187 -4901 138231 -2671
rect 138093 -6543 138108 -4901
rect 138215 -6543 138231 -4901
rect 138093 -10448 138128 -6543
rect 138187 -10448 138231 -6543
rect 138093 -10495 138231 -10448
rect 138332 -10658 138360 -2445
rect 138412 -8688 138448 -2445
rect 138412 -8719 138540 -8688
rect 135144 -10677 138360 -10658
rect 135144 -10721 135416 -10677
rect 138307 -10686 138360 -10677
rect 138412 -9890 138540 -9858
rect 138412 -10686 138448 -9890
rect 138307 -10721 138448 -10686
rect 135144 -10736 138448 -10721
<< via1 >>
rect 93083 26668 94358 26831
rect 89611 26603 89663 26614
rect 89611 26424 89614 26603
rect 89614 26424 89660 26603
rect 89660 26424 89663 26603
rect 89611 26414 89663 26424
rect 92207 26603 92259 26614
rect 92207 26424 92252 26603
rect 92252 26424 92259 26603
rect 92207 26414 92259 26424
rect 95669 26224 95721 26424
rect 90501 25847 91780 26064
rect 88829 25746 89205 25803
rect 90131 25464 90264 25566
rect 92723 25464 92856 25566
rect 93085 25029 94355 25244
rect 89611 24975 89663 24986
rect 89611 24796 89614 24975
rect 89614 24796 89660 24975
rect 89660 24796 89663 24975
rect 89611 24786 89663 24796
rect 92207 24975 92259 24986
rect 92207 24796 92252 24975
rect 92252 24796 92259 24975
rect 92207 24786 92259 24796
rect 95563 24596 95615 24796
rect 90505 24220 91784 24437
rect 88825 24118 89205 24175
rect 90131 23836 90264 23938
rect 92723 23836 92856 23938
rect 93087 23409 94357 23624
rect 89611 23347 89663 23358
rect 89611 23168 89614 23347
rect 89614 23168 89660 23347
rect 89660 23168 89663 23347
rect 89611 23158 89663 23168
rect 92207 23347 92259 23358
rect 92207 23168 92252 23347
rect 92252 23168 92259 23347
rect 92207 23158 92259 23168
rect 95481 22968 95533 23168
rect 90501 22589 91780 22806
rect 88822 22490 89205 22547
rect 90131 22208 90264 22310
rect 92723 22208 92856 22310
rect 93083 21776 94353 21991
rect 89611 21719 89663 21730
rect 89611 21540 89614 21719
rect 89614 21540 89660 21719
rect 89660 21540 89663 21719
rect 89611 21530 89663 21540
rect 92207 21719 92259 21730
rect 92207 21540 92252 21719
rect 92252 21540 92259 21719
rect 92207 21530 92259 21540
rect 95391 21340 95443 21540
rect 90501 20963 91780 21180
rect 88822 20862 89205 20919
rect 90131 20580 90264 20682
rect 92723 20580 92856 20682
rect 93088 20248 94360 20363
rect 95788 20142 95969 21281
rect 95969 20142 96002 21281
rect 96166 23457 96194 25099
rect 96194 23457 96253 25099
rect 96253 23457 96273 25099
rect 138109 23457 138129 25099
rect 138129 23457 138188 25099
rect 138188 23457 138216 25099
rect 138380 20142 138413 21281
rect 138413 20142 138541 21281
rect 89432 10142 89560 11281
rect 89560 10142 89593 11281
rect 89757 13457 89785 15099
rect 89785 13457 89844 15099
rect 89844 13457 89864 15099
rect 138108 13457 138128 15099
rect 138128 13457 138187 15099
rect 138187 13457 138215 15099
rect 138379 10142 138412 11281
rect 138412 10142 138540 11281
rect 89432 142 89560 1281
rect 89560 142 89593 1281
rect 89757 3457 89785 5099
rect 89785 3457 89844 5099
rect 89844 3457 89864 5099
rect 138108 3457 138128 5099
rect 138128 3457 138187 5099
rect 138187 3457 138215 5099
rect 138379 142 138412 1281
rect 138412 142 138540 1281
rect 138108 -6543 138128 -4901
rect 138128 -6543 138187 -4901
rect 138187 -6543 138215 -4901
rect 138379 -9858 138412 -8719
rect 138412 -9858 138540 -8719
<< metal2 >>
rect 89297 28530 103505 28578
rect 88811 26651 89205 26894
rect 88811 25803 88842 26651
rect 89174 25803 89205 26651
rect 88811 25746 88829 25803
rect 88811 25513 88842 25746
rect 89174 25513 89205 25746
rect 88811 24175 89205 25513
rect 88811 24118 88825 24175
rect 88811 22547 89205 24118
rect 89297 22890 89337 28530
rect 89483 28434 103347 28482
rect 89483 24670 89523 28434
rect 89617 28338 101890 28386
rect 89617 26624 89657 28338
rect 89753 28242 101702 28290
rect 89611 26614 89663 26624
rect 89611 26406 89663 26414
rect 89753 25978 89793 28242
rect 91895 28146 100302 28194
rect 89617 25938 89793 25978
rect 90488 26064 91793 26901
rect 89617 24996 89657 25938
rect 90488 25847 90501 26064
rect 91780 25847 91793 26064
rect 90110 25566 90280 25582
rect 90110 25539 90131 25566
rect 89750 25499 90131 25539
rect 89611 24986 89663 24996
rect 89611 24778 89663 24786
rect 89483 24630 89657 24670
rect 89617 23368 89657 24630
rect 89611 23358 89663 23368
rect 89611 23150 89663 23158
rect 89297 22850 89657 22890
rect 88811 22490 88822 22547
rect 88811 20919 89205 22490
rect 89617 21740 89657 22850
rect 89611 21730 89663 21740
rect 89611 21522 89663 21530
rect 88811 20862 88822 20919
rect 88811 20101 89205 20862
rect 89750 19478 89790 25499
rect 90110 25464 90131 25499
rect 90264 25464 90280 25566
rect 90110 25448 90280 25464
rect 90488 25080 91793 25847
rect 90488 24437 90532 25080
rect 91734 24437 91793 25080
rect 90488 24220 90505 24437
rect 91784 24220 91793 24437
rect 90110 23938 90280 23954
rect 90110 23897 90131 23938
rect 89870 23857 90131 23897
rect 89870 19478 89910 23857
rect 90110 23836 90131 23857
rect 90264 23836 90280 23938
rect 90110 23820 90280 23836
rect 90488 23489 90532 24220
rect 91734 23489 91793 24220
rect 90488 22806 91793 23489
rect 91895 22876 91935 28146
rect 92051 28050 100166 28098
rect 92051 24102 92091 28050
rect 92213 27954 98652 28002
rect 92213 26624 92253 27954
rect 92361 27858 98496 27906
rect 92207 26614 92259 26624
rect 92207 26406 92259 26414
rect 92361 25994 92401 27858
rect 97268 27535 97875 27767
rect 98178 27535 98212 27767
rect 98384 27535 98400 27767
rect 97089 27228 97688 27460
rect 97832 27443 98400 27460
rect 98448 27443 98496 27858
rect 97832 27395 98496 27443
rect 98604 27460 98652 27954
rect 98813 27535 98886 27767
rect 99213 27535 99452 27767
rect 99473 27534 100025 27767
rect 98604 27403 99348 27460
rect 97832 27228 98400 27395
rect 98663 27228 99348 27403
rect 99742 27444 99837 27460
rect 100118 27444 100166 28050
rect 99742 27396 100166 27444
rect 100254 27460 100302 28146
rect 100455 27535 100488 27767
rect 100815 27535 101556 27767
rect 99742 27389 99837 27396
rect 99741 27228 99837 27389
rect 100254 27228 100920 27460
rect 101347 27449 101556 27460
rect 101654 27449 101702 28242
rect 101347 27401 101702 27449
rect 101842 27460 101890 28338
rect 102053 27535 102090 27767
rect 102417 27535 103234 27767
rect 101347 27228 101556 27401
rect 101842 27384 102516 27460
rect 101882 27228 102516 27384
rect 102961 27440 103139 27460
rect 103299 27440 103347 28434
rect 102961 27392 103347 27440
rect 103457 27460 103505 28530
rect 103660 27535 103692 27767
rect 104019 27535 105294 27767
rect 105621 27535 106896 27767
rect 107223 27535 108498 27767
rect 108825 27535 113304 27767
rect 113631 27535 119712 27767
rect 120039 27535 120780 27767
rect 121107 27535 122916 27767
rect 123243 27535 130926 27767
rect 131253 27535 137417 27767
rect 102961 27228 103139 27392
rect 103457 27381 137257 27460
rect 103481 27228 137257 27381
rect 97847 27227 97887 27228
rect 100254 27227 100302 27228
rect 92213 25954 92401 25994
rect 93070 26831 94373 26886
rect 93070 26668 93083 26831
rect 94358 26668 94373 26831
rect 96765 26827 137661 27065
rect 92213 24996 92253 25954
rect 92702 25566 92872 25582
rect 92702 25539 92723 25566
rect 92342 25499 92723 25539
rect 92207 24986 92259 24996
rect 92207 24778 92259 24786
rect 92051 24062 92253 24102
rect 92213 23368 92253 24062
rect 92207 23358 92259 23368
rect 92207 23150 92259 23158
rect 91895 22836 92253 22876
rect 90488 22589 90501 22806
rect 91780 22589 91793 22806
rect 90110 22310 90280 22326
rect 90110 22274 90131 22310
rect 89990 22234 90131 22274
rect 89990 19478 90030 22234
rect 90110 22208 90131 22234
rect 90264 22208 90280 22310
rect 90110 22192 90280 22208
rect 90488 21180 91793 22589
rect 92213 21740 92253 22836
rect 92207 21730 92259 21740
rect 92207 21522 92259 21530
rect 90488 20963 90501 21180
rect 91780 20963 91793 21180
rect 90110 20682 90280 20698
rect 90110 20580 90131 20682
rect 90264 20580 90280 20682
rect 90110 20564 90280 20580
rect 90110 19478 90150 20564
rect 90488 20190 91793 20963
rect 92342 19478 92382 25499
rect 92702 25464 92723 25499
rect 92856 25464 92872 25566
rect 92702 25448 92872 25464
rect 93070 25244 94373 26668
rect 96442 26496 96471 26730
rect 96726 26496 96773 26730
rect 137539 26496 137661 26730
rect 137911 26496 137940 26730
rect 95669 26424 95721 26432
rect 95669 26218 95721 26224
rect 94849 26144 94979 26184
rect 93070 25029 93085 25244
rect 94355 25029 94373 25244
rect 92702 23938 92872 23954
rect 92702 23897 92723 23938
rect 92462 23857 92723 23897
rect 92462 19478 92502 23857
rect 92702 23836 92723 23857
rect 92856 23836 92872 23938
rect 92702 23820 92872 23836
rect 93070 23624 94373 25029
rect 95563 24796 95615 24804
rect 95563 24590 95615 24596
rect 93070 23409 93087 23624
rect 94357 23409 94373 23624
rect 92702 22310 92872 22326
rect 92702 22274 92723 22310
rect 92578 22234 92723 22274
rect 92578 19896 92622 22234
rect 92702 22208 92723 22234
rect 92856 22208 92872 22310
rect 92702 22192 92872 22208
rect 93070 21991 94373 23409
rect 95481 23168 95533 23176
rect 95481 22962 95533 22968
rect 93070 21776 93083 21991
rect 94353 21776 94373 21991
rect 93070 21285 94373 21776
rect 95391 21540 95443 21548
rect 95391 21334 95443 21340
rect 92702 20682 92872 20698
rect 92702 20580 92723 20682
rect 92856 20580 92872 20682
rect 92702 20564 92872 20580
rect 92578 19478 92618 19896
rect 92702 19478 92742 20564
rect 93070 20363 93104 21285
rect 94346 20363 94373 21285
rect 93070 20248 93088 20363
rect 94360 20248 94373 20363
rect 93070 20140 93104 20248
rect 94346 20140 94373 20248
rect 93070 20100 94373 20140
rect 95397 19090 95437 21334
rect 95487 19180 95527 22962
rect 95569 19262 95609 24590
rect 95675 19348 95715 26218
rect 96765 25496 137661 25730
rect 137541 25495 137661 25496
rect 96111 25099 96302 25122
rect 96111 23457 96166 25099
rect 96273 23457 96302 25099
rect 138080 25099 138271 25122
rect 96765 24492 137617 24726
rect 96111 23438 96302 23457
rect 96443 23438 96472 23672
rect 96727 23438 96773 23672
rect 137545 23538 137655 23672
rect 137413 23454 137655 23538
rect 137545 23438 137655 23454
rect 137910 23438 137939 23672
rect 138080 23457 138109 25099
rect 138216 23457 138271 25099
rect 138080 23438 138271 23457
rect 126302 23263 137661 23280
rect 137413 23179 137661 23263
rect 137335 23177 137661 23179
rect 126302 23042 137661 23177
rect 96784 22018 137605 22256
rect 95759 21281 96023 21312
rect 95759 20142 95788 21281
rect 96002 20142 96023 21281
rect 138359 21281 138541 21312
rect 95759 20110 96023 20142
rect 96784 20046 137661 20284
rect 138359 20142 138380 21281
rect 138359 20110 138541 20142
rect 97081 19666 97196 19837
rect 97313 19666 97691 19837
rect 98171 19779 98770 19837
rect 97081 19649 97691 19666
rect 98152 19649 98770 19779
rect 99209 19717 99839 19837
rect 99201 19649 99839 19717
rect 100278 19649 100909 19837
rect 101348 19718 137222 19837
rect 101334 19649 137222 19718
rect 97246 19393 97856 19581
rect 98152 19348 98192 19649
rect 98300 19393 98472 19581
rect 98799 19393 98935 19581
rect 95675 19308 98192 19348
rect 99201 19262 99241 19649
rect 99374 19393 99520 19581
rect 99847 19393 99996 19581
rect 95569 19222 99241 19262
rect 100279 19180 100319 19649
rect 100435 19393 100525 19581
rect 100852 19393 101072 19581
rect 95487 19140 100319 19180
rect 101334 19090 101374 19649
rect 132640 19581 132967 19587
rect 101511 19393 101604 19581
rect 101931 19393 137385 19581
rect 95397 19050 101374 19090
rect 130876 18530 138540 18578
rect 90556 17535 92448 17767
rect 92775 17535 103128 17767
rect 103455 17535 111138 17767
rect 111465 17535 113274 17767
rect 113601 17535 114342 17767
rect 114669 17535 120750 17767
rect 121077 17535 125556 17767
rect 125883 17535 127158 17767
rect 127485 17535 128760 17767
rect 129087 17535 130362 17767
rect 130689 17535 130721 17767
rect 130876 17460 130924 18530
rect 90716 17381 130924 17460
rect 131034 18434 138540 18482
rect 131034 17440 131082 18434
rect 132491 18338 138540 18386
rect 131147 17535 131964 17767
rect 132291 17535 132328 17767
rect 132491 17460 132539 18338
rect 131242 17440 131420 17460
rect 131034 17392 131420 17440
rect 90716 17228 130900 17381
rect 131242 17228 131420 17392
rect 131865 17384 132539 17460
rect 132679 18242 138540 18290
rect 132679 17449 132727 18242
rect 134079 18146 138540 18194
rect 132825 17535 133566 17767
rect 133893 17535 133926 17767
rect 134079 17460 134127 18146
rect 132825 17449 133034 17460
rect 132679 17401 133034 17449
rect 131865 17228 132499 17384
rect 132825 17228 133034 17401
rect 133461 17228 134127 17460
rect 134215 18050 138540 18098
rect 134215 17444 134263 18050
rect 135729 17954 138540 18002
rect 134356 17534 134908 17767
rect 134929 17535 135168 17767
rect 135495 17535 135568 17767
rect 135729 17460 135777 17954
rect 134544 17444 134639 17460
rect 134215 17396 134639 17444
rect 134544 17389 134639 17396
rect 135033 17403 135777 17460
rect 135885 17858 138540 17906
rect 135885 17443 135933 17858
rect 135981 17535 135997 17767
rect 136169 17535 136203 17767
rect 136506 17535 137113 17767
rect 135981 17443 136549 17460
rect 134544 17228 134640 17389
rect 135033 17228 135718 17403
rect 135885 17395 136549 17443
rect 135981 17228 136549 17395
rect 136693 17228 137292 17460
rect 134079 17227 134127 17228
rect 136494 17227 136534 17228
rect 90312 16827 137616 17065
rect 90033 16496 90062 16730
rect 90317 16496 90434 16730
rect 137608 16496 137655 16730
rect 137910 16496 137939 16730
rect 90312 15496 137616 15730
rect 90312 15495 90432 15496
rect 89702 15099 89893 15122
rect 89702 13457 89757 15099
rect 89864 13457 89893 15099
rect 138079 15099 138270 15122
rect 90356 14492 137616 14726
rect 89702 13438 89893 13457
rect 90034 13438 90063 13672
rect 90318 13538 90364 13672
rect 90318 13454 90560 13538
rect 90318 13438 90364 13454
rect 137608 13438 137654 13672
rect 137909 13438 137938 13672
rect 138079 13457 138108 15099
rect 138215 13457 138270 15099
rect 138079 13438 138270 13457
rect 90312 13263 108079 13280
rect 90312 13179 90560 13263
rect 90312 13177 90638 13179
rect 90312 13042 108079 13177
rect 90368 12018 137597 12256
rect 89432 11281 89614 11312
rect 89593 10142 89614 11281
rect 138358 11281 138540 11312
rect 89432 10110 89614 10142
rect 90312 10046 137597 10284
rect 138358 10142 138379 11281
rect 138358 10110 138540 10142
rect 90751 9718 133033 9837
rect 90751 9649 133047 9718
rect 133472 9649 134103 9837
rect 134542 9717 135172 9837
rect 135611 9779 136210 9837
rect 134542 9649 135180 9717
rect 135611 9649 136229 9779
rect 136690 9666 137068 9837
rect 137185 9666 137300 9837
rect 136690 9649 137300 9666
rect 101414 9581 101741 9587
rect 90588 9393 132450 9581
rect 132777 9393 132870 9581
rect 133007 9090 133047 9649
rect 133309 9393 133529 9581
rect 133856 9393 133946 9581
rect 134062 9180 134102 9649
rect 134385 9393 134534 9581
rect 134861 9393 135007 9581
rect 135140 9262 135180 9649
rect 135446 9393 135582 9581
rect 135909 9393 136081 9581
rect 136189 9348 136229 9649
rect 136525 9393 137135 9581
rect 136189 9308 138540 9348
rect 135140 9222 138540 9262
rect 134062 9140 138540 9180
rect 133007 9050 138540 9090
rect 130876 8530 138540 8578
rect 90556 7535 92448 7767
rect 92775 7535 103128 7767
rect 103455 7535 111138 7767
rect 111465 7535 113274 7767
rect 113601 7535 114342 7767
rect 114669 7535 120750 7767
rect 121077 7535 125556 7767
rect 125883 7535 127158 7767
rect 127485 7535 128760 7767
rect 129087 7535 130362 7767
rect 130689 7535 130721 7767
rect 130876 7460 130924 8530
rect 90716 7381 130924 7460
rect 131034 8434 138540 8482
rect 131034 7440 131082 8434
rect 132491 8338 138540 8386
rect 131147 7535 131964 7767
rect 132291 7535 132328 7767
rect 132491 7460 132539 8338
rect 131242 7440 131420 7460
rect 131034 7392 131420 7440
rect 90716 7228 130900 7381
rect 131242 7228 131420 7392
rect 131865 7384 132539 7460
rect 132679 8242 138540 8290
rect 132679 7449 132727 8242
rect 134079 8146 138540 8194
rect 132825 7535 133566 7767
rect 133893 7535 133926 7767
rect 134079 7460 134127 8146
rect 132825 7449 133034 7460
rect 132679 7401 133034 7449
rect 131865 7228 132499 7384
rect 132825 7228 133034 7401
rect 133461 7228 134127 7460
rect 134215 8050 138540 8098
rect 134215 7444 134263 8050
rect 135729 7954 138540 8002
rect 134356 7534 134908 7767
rect 134929 7535 135168 7767
rect 135495 7535 135568 7767
rect 135729 7460 135777 7954
rect 134544 7444 134639 7460
rect 134215 7396 134639 7444
rect 134544 7389 134639 7396
rect 135033 7403 135777 7460
rect 135885 7858 138540 7906
rect 135885 7443 135933 7858
rect 135981 7535 135997 7767
rect 136169 7535 136203 7767
rect 136506 7535 137113 7767
rect 135981 7443 136549 7460
rect 134544 7228 134640 7389
rect 135033 7228 135718 7403
rect 135885 7395 136549 7443
rect 135981 7228 136549 7395
rect 136693 7228 137292 7460
rect 134079 7227 134127 7228
rect 136494 7227 136534 7228
rect 90312 6827 137616 7065
rect 90033 6496 90062 6730
rect 90317 6496 90434 6730
rect 137608 6496 137655 6730
rect 137910 6496 137939 6730
rect 90312 5496 137616 5730
rect 90312 5495 90432 5496
rect 89702 5099 89893 5122
rect 89702 3457 89757 5099
rect 89864 3457 89893 5099
rect 138079 5099 138270 5122
rect 90356 4492 137616 4726
rect 89702 3438 89893 3457
rect 90034 3438 90063 3672
rect 90318 3538 90364 3672
rect 90318 3454 90560 3538
rect 90318 3438 90364 3454
rect 137608 3438 137654 3672
rect 137909 3438 137938 3672
rect 138079 3457 138108 5099
rect 138215 3457 138270 5099
rect 138079 3438 138270 3457
rect 90312 3263 108079 3280
rect 90312 3179 90560 3263
rect 90312 3177 90638 3179
rect 90312 3042 108079 3177
rect 90368 2018 137597 2256
rect 89432 1281 89614 1312
rect 89593 142 89614 1281
rect 138358 1281 138540 1312
rect 89432 110 89614 142
rect 90312 46 137597 284
rect 138358 142 138379 1281
rect 138358 110 138540 142
rect 90751 -282 133033 -163
rect 90751 -351 133047 -282
rect 133472 -351 134103 -163
rect 134542 -283 135172 -163
rect 135611 -221 136210 -163
rect 134542 -351 135180 -283
rect 135611 -351 136229 -221
rect 136690 -334 137068 -163
rect 137185 -334 137300 -163
rect 136690 -351 137300 -334
rect 101414 -419 101741 -413
rect 90588 -607 132450 -419
rect 132777 -607 132870 -419
rect 133007 -910 133047 -351
rect 133309 -607 133529 -419
rect 133856 -607 133946 -419
rect 134062 -820 134102 -351
rect 134385 -607 134534 -419
rect 134861 -607 135007 -419
rect 135140 -738 135180 -351
rect 135446 -607 135582 -419
rect 135909 -607 136081 -419
rect 136189 -652 136229 -351
rect 136525 -607 137135 -419
rect 136189 -692 138540 -652
rect 135140 -778 138540 -738
rect 134062 -860 138540 -820
rect 133007 -950 138540 -910
rect 135412 -2465 137704 -2233
rect 135572 -2772 137704 -2540
rect 135168 -3173 137704 -2935
rect 135168 -3504 135290 -3270
rect 137608 -3504 137655 -3270
rect 137910 -3504 137939 -3270
rect 135168 -4504 137704 -4270
rect 135168 -4505 135288 -4504
rect 138079 -4901 138270 -4878
rect 135224 -5508 137704 -5274
rect 137608 -6462 137654 -6328
rect 135215 -6546 135416 -6462
rect 137608 -6562 137654 -6546
rect 137909 -6562 137938 -6328
rect 138079 -6543 138108 -4901
rect 138215 -6543 138270 -4901
rect 138079 -6562 138270 -6543
rect 135168 -6737 137704 -6720
rect 135168 -6821 135416 -6737
rect 135168 -6823 135494 -6821
rect 135168 -6958 137704 -6823
rect 135224 -7982 137704 -7744
rect 138358 -8719 138540 -8688
rect 135168 -9954 137704 -9716
rect 138358 -9858 138379 -8719
rect 138358 -9890 138540 -9858
rect 135607 -10351 137704 -10163
rect 135444 -10607 137704 -10419
<< via2 >>
rect 88842 25803 89174 26651
rect 88842 25746 89174 25803
rect 88842 25513 89174 25746
rect 90532 24437 91734 25080
rect 90532 24220 91734 24437
rect 90532 23489 91734 24220
rect 98212 27535 98384 27767
rect 98886 27535 99213 27767
rect 100488 27535 100815 27767
rect 102090 27535 102417 27767
rect 103692 27535 104019 27767
rect 105294 27535 105621 27767
rect 106896 27535 107223 27767
rect 108498 27535 108825 27767
rect 113304 27535 113631 27767
rect 119712 27535 120039 27767
rect 120780 27535 121107 27767
rect 122916 27535 123243 27767
rect 130926 27535 131253 27767
rect 96471 26496 96726 26730
rect 137661 26496 137911 26730
rect 93104 20363 94346 21285
rect 93104 20248 94346 20363
rect 93104 20140 94346 20248
rect 96166 23457 96273 25099
rect 96472 23438 96727 23672
rect 97235 23454 137413 23538
rect 137655 23438 137910 23672
rect 138109 23457 138216 25099
rect 97234 23179 137413 23263
rect 125319 23177 137335 23179
rect 95788 20142 96002 21281
rect 138380 20142 138541 21281
rect 97196 19666 97313 19837
rect 98472 19393 98799 19581
rect 99520 19393 99847 19581
rect 100525 19393 100852 19581
rect 101604 19393 101931 19581
rect 92448 17535 92775 17767
rect 103128 17535 103455 17767
rect 111138 17535 111465 17767
rect 113274 17535 113601 17767
rect 114342 17535 114669 17767
rect 120750 17535 121077 17767
rect 125556 17535 125883 17767
rect 127158 17535 127485 17767
rect 128760 17535 129087 17767
rect 130362 17535 130689 17767
rect 131964 17535 132291 17767
rect 133566 17535 133893 17767
rect 135168 17535 135495 17767
rect 135997 17535 136169 17767
rect 90062 16496 90317 16730
rect 137655 16496 137910 16730
rect 89757 13457 89864 15099
rect 90063 13438 90318 13672
rect 90560 13454 137146 13538
rect 137654 13438 137909 13672
rect 138108 13457 138215 15099
rect 90560 13179 137147 13263
rect 90638 13177 109062 13179
rect 89432 10142 89593 11281
rect 138379 10142 138540 11281
rect 137068 9666 137185 9837
rect 132450 9393 132777 9581
rect 133529 9393 133856 9581
rect 134534 9393 134861 9581
rect 135582 9393 135909 9581
rect 92448 7535 92775 7767
rect 103128 7535 103455 7767
rect 111138 7535 111465 7767
rect 113274 7535 113601 7767
rect 114342 7535 114669 7767
rect 120750 7535 121077 7767
rect 125556 7535 125883 7767
rect 127158 7535 127485 7767
rect 128760 7535 129087 7767
rect 130362 7535 130689 7767
rect 131964 7535 132291 7767
rect 133566 7535 133893 7767
rect 135168 7535 135495 7767
rect 135997 7535 136169 7767
rect 90062 6496 90317 6730
rect 137655 6496 137910 6730
rect 89757 3457 89864 5099
rect 90063 3438 90318 3672
rect 90560 3454 137146 3538
rect 137654 3438 137909 3672
rect 138108 3457 138215 5099
rect 90560 3179 137147 3263
rect 90638 3177 109062 3179
rect 89432 142 89593 1281
rect 138379 142 138540 1281
rect 137068 -334 137185 -163
rect 132450 -607 132777 -419
rect 133529 -607 133856 -419
rect 134534 -607 134861 -419
rect 135582 -607 135909 -419
rect 137655 -3504 137910 -3270
rect 137654 -6462 137909 -6328
rect 135416 -6546 137909 -6462
rect 137654 -6562 137909 -6546
rect 138108 -6543 138215 -4901
rect 135416 -6821 137704 -6737
rect 135494 -6823 137704 -6821
rect 138379 -9858 138540 -8719
<< metal3 >>
rect 98162 27767 98401 28868
rect 98162 27535 98212 27767
rect 98384 27535 98401 27767
rect 98162 27514 98401 27535
rect 98872 27767 99230 28868
rect 98872 27535 98886 27767
rect 99213 27535 99230 27767
rect 98872 27514 99230 27535
rect 100474 27767 100832 28868
rect 100474 27535 100488 27767
rect 100815 27535 100832 27767
rect 100474 27514 100832 27535
rect 102076 27767 102434 28868
rect 102076 27535 102090 27767
rect 102417 27535 102434 27767
rect 102076 27514 102434 27535
rect 103678 27767 104036 28868
rect 103678 27535 103692 27767
rect 104019 27535 104036 27767
rect 103678 27514 104036 27535
rect 105280 27767 105638 28868
rect 105280 27535 105294 27767
rect 105621 27535 105638 27767
rect 105280 27514 105638 27535
rect 106882 27767 107240 28868
rect 106882 27535 106896 27767
rect 107223 27535 107240 27767
rect 106882 27514 107240 27535
rect 108484 27767 108842 28868
rect 108484 27535 108498 27767
rect 108825 27535 108842 27767
rect 108484 27469 108842 27535
rect 113290 27767 113648 28868
rect 113290 27535 113304 27767
rect 113631 27535 113648 27767
rect 113290 27514 113648 27535
rect 119698 27767 120056 28868
rect 119698 27535 119712 27767
rect 120039 27535 120056 27767
rect 119698 27514 120056 27535
rect 120766 27767 121124 28868
rect 120766 27535 120780 27767
rect 121107 27535 121124 27767
rect 120766 27514 121124 27535
rect 122902 27767 123260 28868
rect 130912 28236 131270 28868
rect 130911 27900 131271 28236
rect 122902 27535 122916 27767
rect 123243 27535 123260 27767
rect 122902 27514 123260 27535
rect 130912 27767 131270 27900
rect 130912 27535 130926 27767
rect 131253 27535 131270 27767
rect 130912 27514 131270 27535
rect 96461 26730 96739 26767
rect 88812 26651 89205 26686
rect 88812 25513 88842 26651
rect 89174 25513 89205 26651
rect 88812 25484 89205 25513
rect 96461 26496 96471 26730
rect 96726 26496 96739 26730
rect 90487 25080 91793 25123
rect 90487 23489 90532 25080
rect 91734 23489 91793 25080
rect 90487 23436 91793 23489
rect 96133 25099 96302 25121
rect 96133 23457 96166 25099
rect 96273 23457 96302 25099
rect 96133 23438 96302 23457
rect 96461 23672 96739 26496
rect 137643 26730 137921 26767
rect 137643 26496 137661 26730
rect 137911 26496 137921 26730
rect 137643 23672 137921 26496
rect 96461 23438 96472 23672
rect 96727 23627 137655 23672
rect 96727 23453 97234 23627
rect 137413 23453 137655 23627
rect 96727 23438 137655 23453
rect 137910 23438 137921 23672
rect 138080 25099 138249 25121
rect 138080 23457 138109 25099
rect 138216 23457 138249 25099
rect 138080 23438 138249 23457
rect 93072 21285 94372 21313
rect 93072 20140 93104 21285
rect 94346 20140 94372 21285
rect 93072 20113 94372 20140
rect 95759 21281 96023 21312
rect 95759 20142 95788 21281
rect 96002 20142 96023 21281
rect 95759 20110 96023 20142
rect 96461 20054 96739 23438
rect 96842 23264 137538 23280
rect 96842 23090 97234 23264
rect 137413 23090 137538 23264
rect 96842 23088 125319 23090
rect 137335 23088 137538 23090
rect 96842 23042 137538 23088
rect 137643 20054 137921 23438
rect 138359 21281 138547 21312
rect 138359 20142 138380 21281
rect 138541 20142 138547 21281
rect 138359 20110 138547 20142
rect 97187 19837 97321 19853
rect 97187 19666 97196 19837
rect 97313 19666 97321 19837
rect 97187 19661 97321 19666
rect 98454 19581 98816 19603
rect 98454 19578 98472 19581
rect 98449 19393 98472 19578
rect 98799 19393 98816 19581
rect 98449 19284 98816 19393
rect 99502 19581 99864 19603
rect 99502 19393 99520 19581
rect 99847 19393 99864 19581
rect 99502 19284 99864 19393
rect 100507 19581 100869 19603
rect 100507 19393 100525 19581
rect 100852 19393 100869 19581
rect 100507 19284 100869 19393
rect 101586 19581 101948 19603
rect 101586 19393 101604 19581
rect 101931 19393 101948 19581
rect 101586 19284 101948 19393
rect 92431 17767 92789 18868
rect 103111 18236 103469 18868
rect 103110 17900 103470 18236
rect 92431 17535 92448 17767
rect 92775 17535 92789 17767
rect 92431 17514 92789 17535
rect 103111 17767 103469 17900
rect 103111 17535 103128 17767
rect 103455 17535 103469 17767
rect 103111 17514 103469 17535
rect 111121 17767 111479 18868
rect 111121 17535 111138 17767
rect 111465 17535 111479 17767
rect 111121 17514 111479 17535
rect 113257 17767 113615 18868
rect 113257 17535 113274 17767
rect 113601 17535 113615 17767
rect 113257 17514 113615 17535
rect 114325 17767 114683 18868
rect 114325 17535 114342 17767
rect 114669 17535 114683 17767
rect 114325 17514 114683 17535
rect 120733 17767 121091 18868
rect 120733 17535 120750 17767
rect 121077 17535 121091 17767
rect 120733 17514 121091 17535
rect 125539 17767 125897 18868
rect 125539 17535 125556 17767
rect 125883 17535 125897 17767
rect 125539 17469 125897 17535
rect 127141 17767 127499 18868
rect 127141 17535 127158 17767
rect 127485 17535 127499 17767
rect 127141 17514 127499 17535
rect 128743 17767 129101 18868
rect 128743 17535 128760 17767
rect 129087 17535 129101 17767
rect 128743 17514 129101 17535
rect 130345 17767 130703 18868
rect 130345 17535 130362 17767
rect 130689 17535 130703 17767
rect 130345 17514 130703 17535
rect 131947 17767 132305 18868
rect 131947 17535 131964 17767
rect 132291 17535 132305 17767
rect 131947 17514 132305 17535
rect 133549 17767 133907 18868
rect 133549 17535 133566 17767
rect 133893 17535 133907 17767
rect 133549 17514 133907 17535
rect 135151 17767 135509 18868
rect 135151 17535 135168 17767
rect 135495 17535 135509 17767
rect 135151 17514 135509 17535
rect 135980 17767 136219 18868
rect 135980 17535 135997 17767
rect 136169 17535 136219 17767
rect 135980 17514 136219 17535
rect 90052 16730 90330 16767
rect 90052 16496 90062 16730
rect 90317 16496 90330 16730
rect 89724 15099 89893 15121
rect 89724 13457 89757 15099
rect 89864 13457 89893 15099
rect 89724 13438 89893 13457
rect 90052 13672 90330 16496
rect 137642 16730 137920 16767
rect 137642 16496 137655 16730
rect 137910 16496 137920 16730
rect 137642 13672 137920 16496
rect 90052 13438 90063 13672
rect 90318 13627 137654 13672
rect 90318 13453 90560 13627
rect 137147 13453 137654 13627
rect 90318 13438 137654 13453
rect 137909 13438 137920 13672
rect 138079 15099 138248 15121
rect 138079 13457 138108 15099
rect 138215 13457 138248 15099
rect 138079 13438 138248 13457
rect 89427 11281 89614 11312
rect 89427 10142 89432 11281
rect 89593 10142 89614 11281
rect 89427 10110 89614 10142
rect 90052 10054 90330 13438
rect 90406 13264 137539 13280
rect 90406 13090 90560 13264
rect 137147 13090 137539 13264
rect 90406 13088 90638 13090
rect 109062 13088 137539 13090
rect 90406 13042 137539 13088
rect 137642 10054 137920 13438
rect 138358 11281 138545 11312
rect 138358 10142 138379 11281
rect 138540 10142 138545 11281
rect 138358 10110 138545 10142
rect 137060 9837 137194 9853
rect 137060 9666 137068 9837
rect 137185 9666 137194 9837
rect 137060 9661 137194 9666
rect 132433 9581 132795 9603
rect 132433 9393 132450 9581
rect 132777 9393 132795 9581
rect 132433 9284 132795 9393
rect 133512 9581 133874 9603
rect 133512 9393 133529 9581
rect 133856 9393 133874 9581
rect 133512 9284 133874 9393
rect 134517 9581 134879 9603
rect 134517 9393 134534 9581
rect 134861 9393 134879 9581
rect 134517 9284 134879 9393
rect 135565 9581 135927 9603
rect 135565 9393 135582 9581
rect 135909 9578 135927 9581
rect 135909 9393 135932 9578
rect 135565 9284 135932 9393
rect 92431 7767 92789 8868
rect 103111 8236 103469 8868
rect 103110 7900 103470 8236
rect 92431 7535 92448 7767
rect 92775 7535 92789 7767
rect 92431 7514 92789 7535
rect 103111 7767 103469 7900
rect 103111 7535 103128 7767
rect 103455 7535 103469 7767
rect 103111 7514 103469 7535
rect 111121 7767 111479 8868
rect 111121 7535 111138 7767
rect 111465 7535 111479 7767
rect 111121 7514 111479 7535
rect 113257 7767 113615 8868
rect 113257 7535 113274 7767
rect 113601 7535 113615 7767
rect 113257 7514 113615 7535
rect 114325 7767 114683 8868
rect 114325 7535 114342 7767
rect 114669 7535 114683 7767
rect 114325 7514 114683 7535
rect 120733 7767 121091 8868
rect 120733 7535 120750 7767
rect 121077 7535 121091 7767
rect 120733 7514 121091 7535
rect 125539 7767 125897 8868
rect 125539 7535 125556 7767
rect 125883 7535 125897 7767
rect 125539 7469 125897 7535
rect 127141 7767 127499 8868
rect 127141 7535 127158 7767
rect 127485 7535 127499 7767
rect 127141 7514 127499 7535
rect 128743 7767 129101 8868
rect 128743 7535 128760 7767
rect 129087 7535 129101 7767
rect 128743 7514 129101 7535
rect 130345 7767 130703 8868
rect 130345 7535 130362 7767
rect 130689 7535 130703 7767
rect 130345 7514 130703 7535
rect 131947 7767 132305 8868
rect 131947 7535 131964 7767
rect 132291 7535 132305 7767
rect 131947 7514 132305 7535
rect 133549 7767 133907 8868
rect 133549 7535 133566 7767
rect 133893 7535 133907 7767
rect 133549 7514 133907 7535
rect 135151 7767 135509 8868
rect 135151 7535 135168 7767
rect 135495 7535 135509 7767
rect 135151 7514 135509 7535
rect 135980 7767 136219 8868
rect 135980 7535 135997 7767
rect 136169 7535 136219 7767
rect 135980 7514 136219 7535
rect 90052 6730 90330 6767
rect 90052 6496 90062 6730
rect 90317 6496 90330 6730
rect 89724 5099 89893 5121
rect 89724 3457 89757 5099
rect 89864 3457 89893 5099
rect 89724 3438 89893 3457
rect 90052 3672 90330 6496
rect 137642 6730 137920 6767
rect 137642 6496 137655 6730
rect 137910 6496 137920 6730
rect 137642 3672 137920 6496
rect 90052 3438 90063 3672
rect 90318 3627 137654 3672
rect 90318 3453 90560 3627
rect 137147 3453 137654 3627
rect 90318 3438 137654 3453
rect 137909 3438 137920 3672
rect 138079 5099 138248 5121
rect 138079 3457 138108 5099
rect 138215 3457 138248 5099
rect 138079 3438 138248 3457
rect 89427 1281 89614 1312
rect 89427 142 89432 1281
rect 89593 142 89614 1281
rect 89427 110 89614 142
rect 90052 54 90330 3438
rect 90417 3264 137539 3280
rect 90417 3090 90560 3264
rect 137147 3090 137539 3264
rect 90417 3088 90638 3090
rect 109062 3088 137539 3090
rect 90417 3042 137539 3088
rect 137642 54 137920 3438
rect 138358 1281 138545 1312
rect 138358 142 138379 1281
rect 138540 142 138545 1281
rect 138358 110 138545 142
rect 137060 -163 137194 -147
rect 137060 -334 137068 -163
rect 137185 -334 137194 -163
rect 137060 -339 137194 -334
rect 132433 -419 132795 -397
rect 132433 -607 132450 -419
rect 132777 -607 132795 -419
rect 132433 -716 132795 -607
rect 133512 -419 133874 -397
rect 133512 -607 133529 -419
rect 133856 -607 133874 -419
rect 133512 -716 133874 -607
rect 134517 -419 134879 -397
rect 134517 -607 134534 -419
rect 134861 -607 134879 -419
rect 134517 -716 134879 -607
rect 135565 -419 135927 -397
rect 135565 -607 135582 -419
rect 135909 -422 135927 -419
rect 135909 -607 135932 -422
rect 135565 -716 135932 -607
rect 137642 -3270 137920 -3233
rect 137642 -3504 137655 -3270
rect 137910 -3504 137920 -3270
rect 137642 -6328 137920 -3504
rect 135208 -6373 137654 -6328
rect 135208 -6547 135416 -6373
rect 135208 -6562 137654 -6547
rect 137909 -6562 137920 -6328
rect 138079 -4901 138248 -4879
rect 138079 -6543 138108 -4901
rect 138215 -6543 138248 -4901
rect 138079 -6562 138248 -6543
rect 137642 -6720 137920 -6562
rect 135219 -6736 137920 -6720
rect 135219 -6910 135416 -6736
rect 135219 -6912 135494 -6910
rect 137704 -6912 137920 -6736
rect 135219 -6958 137920 -6912
rect 137642 -9946 137920 -6958
rect 138358 -8719 138545 -8688
rect 138358 -9858 138379 -8719
rect 138540 -9858 138545 -8719
rect 138358 -9890 138545 -9858
<< via3 >>
rect 88842 25513 89174 26651
rect 90532 23489 91734 25080
rect 96166 23457 96273 25099
rect 97234 23538 137413 23627
rect 97234 23454 97235 23538
rect 97235 23454 137413 23538
rect 97234 23453 137413 23454
rect 138109 23457 138216 25099
rect 93104 20140 94346 21285
rect 95788 20142 96002 21281
rect 97234 23263 137413 23264
rect 97234 23179 137413 23263
rect 97234 23177 125319 23179
rect 125319 23177 137335 23179
rect 137335 23177 137413 23179
rect 97234 23090 137413 23177
rect 125319 23088 137335 23090
rect 138380 20142 138541 21281
rect 89757 13457 89864 15099
rect 90560 13538 137147 13627
rect 90560 13454 137146 13538
rect 137146 13454 137147 13538
rect 90560 13453 137147 13454
rect 138108 13457 138215 15099
rect 89432 10142 89593 11281
rect 90560 13263 137147 13264
rect 90560 13179 137147 13263
rect 90560 13177 90638 13179
rect 90638 13177 109062 13179
rect 109062 13177 137147 13179
rect 90560 13090 137147 13177
rect 90638 13088 109062 13090
rect 138379 10142 138540 11281
rect 89757 3457 89864 5099
rect 90560 3538 137147 3627
rect 90560 3454 137146 3538
rect 137146 3454 137147 3538
rect 90560 3453 137147 3454
rect 138108 3457 138215 5099
rect 89432 142 89593 1281
rect 90560 3263 137147 3264
rect 90560 3179 137147 3263
rect 90560 3177 90638 3179
rect 90638 3177 109062 3179
rect 109062 3177 137147 3179
rect 90560 3090 137147 3177
rect 90638 3088 109062 3090
rect 138379 142 138540 1281
rect 135416 -6462 137654 -6373
rect 137654 -6462 137704 -6373
rect 135416 -6546 137704 -6462
rect 135416 -6547 137654 -6546
rect 137654 -6547 137704 -6546
rect 138108 -6543 138215 -4901
rect 135416 -6737 137704 -6736
rect 135416 -6821 137704 -6737
rect 135416 -6823 135494 -6821
rect 135494 -6823 137704 -6821
rect 135416 -6910 137704 -6823
rect 135494 -6912 137704 -6910
rect 138379 -9858 138540 -8719
<< metal4 >>
rect 88136 26651 96025 26683
rect 88136 25513 88842 26651
rect 89174 25513 96025 26651
rect 88136 25483 96025 25513
rect 138357 25483 138541 26683
rect 88136 25099 138541 25120
rect 88136 25080 96166 25099
rect 88136 23489 90532 25080
rect 91734 23489 96166 25080
rect 88136 23457 96166 23489
rect 96273 23627 138109 25099
rect 96273 23457 97234 23627
rect 88136 23453 97234 23457
rect 137413 23457 138109 23627
rect 138216 23457 138541 25099
rect 137413 23453 138541 23457
rect 88136 23435 138541 23453
rect 88136 23264 138541 23284
rect 88136 23090 97234 23264
rect 137413 23090 138541 23264
rect 88136 23088 125319 23090
rect 137335 23088 138541 23090
rect 88136 21599 138541 23088
rect 88136 21285 96025 21311
rect 88136 20140 93104 21285
rect 94346 21281 96025 21285
rect 94346 20142 95788 21281
rect 96002 20142 96025 21281
rect 94346 20140 96025 20142
rect 88136 20111 96025 20140
rect 138357 21281 138545 21311
rect 138357 20142 138380 21281
rect 138541 20142 138545 21281
rect 138357 20111 138545 20142
rect 89432 15483 89616 16683
rect 138356 15483 138540 16683
rect 89432 15099 138540 15120
rect 89432 13457 89757 15099
rect 89864 13627 138108 15099
rect 89864 13457 90560 13627
rect 89432 13453 90560 13457
rect 137147 13457 138108 13627
rect 138215 13457 138540 15099
rect 137147 13453 138540 13457
rect 89432 13435 138540 13453
rect 89432 13264 138540 13284
rect 89432 13090 90560 13264
rect 137147 13090 138540 13264
rect 89432 13088 90638 13090
rect 109062 13088 138540 13090
rect 89432 11599 138540 13088
rect 89429 11281 89616 11311
rect 89429 10142 89432 11281
rect 89593 10142 89616 11281
rect 89429 10111 89616 10142
rect 138356 11281 138544 11311
rect 138356 10142 138379 11281
rect 138540 10142 138544 11281
rect 138356 10111 138544 10142
rect 89432 5483 89616 6683
rect 138356 5483 138540 6683
rect 89432 5099 138540 5120
rect 89432 3457 89757 5099
rect 89864 3627 138108 5099
rect 89864 3457 90560 3627
rect 89432 3453 90560 3457
rect 137147 3457 138108 3627
rect 138215 3457 138540 5099
rect 137147 3453 138540 3457
rect 89432 3435 138540 3453
rect 89432 3264 138540 3284
rect 89432 3090 90560 3264
rect 137147 3090 138540 3264
rect 89432 3088 90638 3090
rect 109062 3088 138540 3090
rect 89432 1599 138540 3088
rect 89429 1281 89616 1311
rect 89429 142 89432 1281
rect 89593 142 89616 1281
rect 89429 111 89616 142
rect 138356 1281 138543 1311
rect 138356 142 138379 1281
rect 138540 142 138543 1281
rect 138356 111 138543 142
rect 138356 -4517 138540 -3317
rect 135167 -4901 138540 -4880
rect 135167 -6373 138108 -4901
rect 135167 -6547 135416 -6373
rect 137704 -6543 138108 -6373
rect 138215 -6543 138540 -4901
rect 137704 -6547 138540 -6543
rect 135167 -6565 138540 -6547
rect 135168 -6736 138540 -6716
rect 135168 -6910 135416 -6736
rect 135168 -6912 135494 -6910
rect 137704 -6912 138540 -6736
rect 135168 -8401 138540 -6912
rect 138356 -8719 138546 -8689
rect 138356 -9858 138379 -8719
rect 138540 -9858 138546 -8719
rect 138356 -9889 138546 -9858
use bias_nstack  bias_nstack_0
array 0 75 -534 0 0 -4355
timestamp 1717035242
transform 1 0 133578 0 -1 20420
box 3258 -2860 3926 1035
use bias_nstack  bias_nstack_1
array 0 87 -534 0 0 -4355
timestamp 1717035242
transform -1 0 94395 0 -1 10420
box 3258 -2860 3926 1035
use bias_nstack  bias_nstack_2
array 0 87 -534 0 0 -4355
timestamp 1717035242
transform -1 0 94395 0 -1 420
box 3258 -2860 3926 1035
use bias_nstack  bias_nstack_3
array 0 3 -534 0 0 -4355
timestamp 1717035242
transform -1 0 139251 0 -1 -9580
box 3258 -2860 3926 1035
use bias_pstack  bias_pstack_0
array 0 75 534 0 0 -4355
timestamp 1717035242
transform -1 0 139531 0 -1 23826
box 1986 -3967 2714 388
use bias_pstack  bias_pstack_1
array 0 87 534 0 0 -4355
timestamp 1717035242
transform 1 0 88442 0 -1 13826
box 1986 -3967 2714 388
use bias_pstack  bias_pstack_2
array 0 87 534 0 0 -4355
timestamp 1717035242
transform 1 0 88442 0 -1 3826
box 1986 -3967 2714 388
use bias_pstack  bias_pstack_3
array 0 3 534 0 0 -4355
timestamp 1717035242
transform 1 0 133298 0 -1 -6174
box 1986 -3967 2714 388
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform 1 0 94485 0 -1 23514
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_1
timestamp 1715205430
transform 1 0 94485 0 -1 26770
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_8
timestamp 1715205430
transform 1 0 91893 0 1 20258
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_9
timestamp 1715205430
transform 1 0 91893 0 1 23514
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_10
timestamp 1715205430
transform 1 0 91893 0 1 21886
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_11
timestamp 1715205430
transform 1 0 94485 0 1 20258
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_12
timestamp 1715205430
transform 1 0 91893 0 1 25142
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_13
timestamp 1715205430
transform 1 0 94485 0 1 25142
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_14
timestamp 1715205430
transform 1 0 94485 0 -1 21886
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_16
timestamp 1715205430
transform 1 0 94485 0 1 23514
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_17
timestamp 1715205430
transform 1 0 94485 0 1 21886
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_18
timestamp 1715205430
transform 1 0 94485 0 -1 25142
box -66 -43 450 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_8 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform 1 0 92277 0 1 20258
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_9
timestamp 1715205430
transform 1 0 92277 0 1 23514
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_10
timestamp 1715205430
transform 1 0 92277 0 1 21886
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_11
timestamp 1715205430
transform 1 0 94869 0 1 20258
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_12
timestamp 1715205430
transform 1 0 92277 0 1 25142
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_13
timestamp 1715205430
transform 1 0 94869 0 1 25142
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_14
timestamp 1715205430
transform 1 0 94869 0 -1 21886
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_15
timestamp 1715205430
transform 1 0 94869 0 -1 23514
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_16
timestamp 1715205430
transform 1 0 94869 0 1 23514
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_17
timestamp 1715205430
transform 1 0 94869 0 1 21886
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_18
timestamp 1715205430
transform 1 0 94869 0 -1 25142
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_19
timestamp 1715205430
transform 1 0 94869 0 -1 26770
box -66 -43 162 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform 1 0 91893 0 -1 21886
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_7
timestamp 1715205430
transform 1 0 91893 0 -1 23514
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_10
timestamp 1715205430
transform 1 0 91893 0 -1 26770
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_11
timestamp 1715205430
transform 1 0 91893 0 -1 25142
box -66 -43 546 897
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
array 0 1 -2592 0 3 1628
timestamp 1715205430
transform 1 0 92373 0 1 20258
box -66 -43 2178 1671
<< labels >>
flabel metal4 135168 -8401 135401 -6716 0 FreeSans 1600 90 0 0 avss
port 2 nsew
flabel metal4 135167 -6565 135400 -4880 0 FreeSans 1600 90 0 0 avdd
port 1 nsew
flabel metal3 92431 8625 92789 8865 0 FreeSans 1600 90 0 0 idac_src_1000
port 38 nsew
flabel metal3 103111 8625 103469 8865 0 FreeSans 1600 90 0 0 hsxo_src_1000
port 37 nsew
flabel metal3 111121 8625 111479 8865 0 FreeSans 1600 90 0 0 test_src_500
port 36 nsew
flabel metal3 113257 8625 113615 8865 0 FreeSans 1600 90 0 0 user_src_150
port 35 nsew
flabel metal3 114325 8625 114683 8865 0 FreeSans 1600 90 0 0 user_src_50
port 34 nsew
flabel metal3 120733 8625 121091 8865 0 FreeSans 1600 90 0 0 ov_src_600
port 33 nsew
flabel metal3 127141 8625 127499 8865 0 FreeSans 1600 90 0 0 instr2_src_100
port 31 nsew
flabel metal3 128743 8625 129101 8865 0 FreeSans 1600 90 0 0 instr1_src_100
port 30 nsew
flabel metal3 130345 8625 130703 8865 0 FreeSans 1600 90 0 0 hgbw2_src_100
port 29 nsew
flabel metal3 131947 8625 132305 8865 0 FreeSans 1600 90 0 0 hgbw1_src_100
port 28 nsew
flabel metal3 133549 8625 133907 8865 0 FreeSans 1600 90 0 0 lp2_src_100
port 27 nsew
flabel metal3 135151 8625 135509 8865 0 FreeSans 1600 90 0 0 lp1_src_100
port 8 nsew
flabel metal3 135980 8625 136219 8865 0 FreeSans 1600 90 0 0 lsxo_src_50
port 7 nsew
flabel metal3 125539 8625 125897 8865 0 FreeSans 1600 90 0 0 en_comp_trim_n
port 32 nsew
flabel metal4 90311 3435 90544 5120 0 FreeSans 1600 90 0 0 avdd
port 1 nsew
flabel metal4 90312 1599 90545 3284 0 FreeSans 1600 90 0 0 avss
port 2 nsew
flabel metal3 92431 18625 92789 18865 0 FreeSans 1600 90 0 0 idac_src_1000
port 38 nsew
flabel metal3 103111 18625 103469 18865 0 FreeSans 1600 90 0 0 hsxo_src_1000
port 37 nsew
flabel metal3 111121 18625 111479 18865 0 FreeSans 1600 90 0 0 test_src_500
port 36 nsew
flabel metal3 113257 18625 113615 18865 0 FreeSans 1600 90 0 0 user_src_150
port 35 nsew
flabel metal3 114325 18625 114683 18865 0 FreeSans 1600 90 0 0 user_src_50
port 34 nsew
flabel metal3 120733 18625 121091 18865 0 FreeSans 1600 90 0 0 ov_src_600
port 33 nsew
flabel metal3 127141 18625 127499 18865 0 FreeSans 1600 90 0 0 instr2_src_100
port 31 nsew
flabel metal3 128743 18625 129101 18865 0 FreeSans 1600 90 0 0 instr1_src_100
port 30 nsew
flabel metal3 130345 18625 130703 18865 0 FreeSans 1600 90 0 0 hgbw2_src_100
port 29 nsew
flabel metal3 131947 18625 132305 18865 0 FreeSans 1600 90 0 0 hgbw1_src_100
port 28 nsew
flabel metal3 133549 18625 133907 18865 0 FreeSans 1600 90 0 0 lp2_src_100
port 27 nsew
flabel metal3 135151 18625 135509 18865 0 FreeSans 1600 90 0 0 lp1_src_100
port 8 nsew
flabel metal3 135980 18625 136219 18865 0 FreeSans 1600 90 0 0 lsxo_src_50
port 7 nsew
flabel metal3 125539 18625 125897 18865 0 FreeSans 1600 90 0 0 en_comp_trim_n
port 32 nsew
flabel metal4 90311 13435 90544 15120 0 FreeSans 1600 90 0 0 avdd
port 1 nsew
flabel metal4 90312 11599 90545 13284 0 FreeSans 1600 90 0 0 avss
port 2 nsew
flabel metal4 137603 23435 137662 25120 0 FreeSans 1600 90 0 0 avdd
port 1 nsew
flabel metal4 137603 21599 137661 23284 0 FreeSans 1600 90 0 0 avss
port 2 nsew
flabel metal3 108484 28625 108842 28865 0 FreeSans 1600 90 0 0 en_comp_trim_n
port 32 nsew
flabel metal3 98162 28625 98401 28865 0 FreeSans 1600 90 0 0 lsxo_src_50
port 7 nsew
flabel metal3 98872 28625 99230 28865 0 FreeSans 1600 90 0 0 lp1_src_100
port 8 nsew
flabel metal3 100474 28625 100832 28865 0 FreeSans 1600 90 0 0 lp2_src_100
port 27 nsew
flabel metal3 102076 28625 102434 28865 0 FreeSans 1600 90 0 0 hgbw1_src_100
port 28 nsew
flabel metal3 103678 28625 104036 28865 0 FreeSans 1600 90 0 0 hgbw2_src_100
port 29 nsew
flabel metal3 105280 28625 105638 28865 0 FreeSans 1600 90 0 0 instr1_src_100
port 30 nsew
flabel metal3 106882 28625 107240 28865 0 FreeSans 1600 90 0 0 instr2_src_100
port 31 nsew
flabel metal3 113290 28625 113648 28865 0 FreeSans 1600 90 0 0 ov_src_600
port 33 nsew
flabel metal3 119698 28625 120056 28865 0 FreeSans 1600 90 0 0 user_src_50
port 34 nsew
flabel metal3 120766 28625 121124 28865 0 FreeSans 1600 90 0 0 user_src_150
port 35 nsew
flabel metal3 122902 28625 123260 28865 0 FreeSans 1600 90 0 0 test_src_500
port 36 nsew
flabel metal3 130912 28625 131270 28865 0 FreeSans 1600 90 0 0 hsxo_src_1000
port 37 nsew
flabel metal4 88136 25483 88736 26683 0 FreeSans 3200 90 0 0 dvdd
port 3 nsew
flabel metal4 88136 23435 88736 25120 0 FreeSans 3200 90 0 0 avdd
port 1 nsew
flabel metal4 88136 21599 88736 23284 0 FreeSans 3200 90 0 0 avss
port 2 nsew
flabel metal4 88136 20111 88736 21311 0 FreeSans 3200 90 0 0 dvss
port 4 nsew
flabel metal2 92702 19478 92742 19878 0 FreeSans 400 90 0 0 en_snk_test
port 26 nsew
flabel metal2 92578 19478 92618 19853 0 FreeSans 400 90 0 0 en_user2_trim_n
port 16 nsew
flabel metal2 92462 19478 92502 19853 0 FreeSans 400 90 0 0 en_comp_trim_n
port 24 nsew
flabel metal2 92342 19478 92382 19853 0 FreeSans 400 90 0 0 en_hsxo_trim_n
port 25 nsew
flabel metal2 90110 19478 90150 19853 0 FreeSans 400 90 0 0 en_lp2_bias
port 20 nsew
flabel metal2 89990 19478 90030 19853 0 FreeSans 400 90 0 0 en_lp1_trim_p
port 21 nsew
flabel metal2 89870 19478 89910 19853 0 FreeSans 400 90 0 0 en_lsxo_bias
port 23 nsew
flabel metal2 89750 19478 89790 19853 0 FreeSans 400 90 0 0 en_lp1_bias
port 22 nsew
<< end >>
