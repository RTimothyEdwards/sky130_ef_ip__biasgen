magic
tech sky130A
magscale 1 2
timestamp 1720038234
<< viali >>
rect 1082 218 1148 1710
<< metal1 >>
rect 435 7250 5527 7371
rect 856 4999 1685 5067
rect 1078 3439 1162 3440
rect 852 3371 1685 3439
rect 1037 1743 1685 1811
rect 1052 1710 1176 1743
rect 1052 218 1082 1710
rect 1148 218 1176 1710
rect 1052 183 1176 218
rect 1037 115 1685 183
<< metal2 >>
rect 142 34487 182 34862
rect 262 34487 302 34862
rect 382 34487 422 34862
rect 502 34487 542 34862
rect 2734 34487 2774 34862
rect 2854 34487 2894 34862
rect 2970 34487 3010 34862
rect 3094 34462 3134 34862
rect 48508 26791 49914 26810
rect 48508 25622 48529 26791
rect 48833 25622 49574 26791
rect 48508 25616 49574 25622
rect 49888 25616 49914 26791
rect 48508 25597 49914 25616
rect 47968 10123 48017 10357
rect 48511 8284 49913 8311
rect 48511 8280 49576 8284
rect 47877 7213 48035 7273
rect 48511 7160 48546 8280
rect 48816 7160 49576 8280
rect 48511 7150 49576 7160
rect 49888 7150 49913 8284
rect 48511 7127 49913 7150
rect 48035 5092 48038 5326
rect 48035 4088 48038 4322
rect 48035 1614 48047 1852
<< via2 >>
rect 7681 34828 47745 34890
rect 7699 26652 47763 26714
rect 1005 25695 47470 25757
rect 48529 25622 48833 26791
rect 49574 25616 49888 26791
rect 1553 17526 41617 17588
rect 1028 16343 41092 16405
rect 1005 8161 47469 8223
rect 45880 7213 47877 7273
rect 48546 7160 48816 8280
rect 49576 7150 49888 8284
rect 45884 -946 48005 -888
<< metal3 >>
rect 49073 34950 49433 35112
rect 7638 34890 49433 34950
rect 7638 34828 7681 34890
rect 47745 34828 49433 34890
rect 7638 34758 49433 34828
rect 0 34198 246 34232
rect 0 33050 30 34198
rect 220 33050 246 34198
rect 0 33026 246 33050
rect -352 27080 -212 28868
rect -1110 26940 -212 27080
rect -1110 7594 -970 26940
rect 48 26880 188 33026
rect -910 26740 188 26880
rect 7648 26791 48859 26812
rect -910 19396 -770 26740
rect 7648 26714 48529 26791
rect 7648 26652 7699 26714
rect 47763 26652 48529 26714
rect 7648 26576 48529 26652
rect 47807 25858 48529 26576
rect 951 25757 48529 25858
rect 951 25695 1005 25757
rect 47470 25695 48529 25757
rect 951 25622 48529 25695
rect 48833 25622 48859 26791
rect 951 25597 48859 25622
rect -910 19136 8 19396
rect -910 18494 -758 19136
rect -278 18494 8 19136
rect -910 18184 8 18494
rect -910 15748 -770 18184
rect 49073 17659 49433 34758
rect 1478 17588 49433 17659
rect 1478 17526 1553 17588
rect 41617 17526 49433 17588
rect 1478 17464 49433 17526
rect 47867 16464 49433 17464
rect 978 16405 49433 16464
rect 978 16343 1028 16405
rect 41092 16343 49433 16405
rect 978 16269 49433 16343
rect -910 15452 12 15748
rect -910 14810 -756 15452
rect -276 14810 12 15452
rect -910 14536 12 14810
rect -910 7794 -770 14536
rect 960 8280 48855 8312
rect 960 8223 48546 8280
rect 960 8161 1005 8223
rect 47469 8161 48546 8223
rect 960 8087 48546 8161
rect -910 7654 1690 7794
rect -1110 7454 1290 7594
rect 1150 6316 1290 7454
rect 1116 6296 1370 6316
rect 1116 4936 1132 6296
rect 1344 4936 1370 6296
rect 1116 4920 1370 4936
rect 1550 296 1690 7654
rect 47877 7363 48546 8087
rect 45838 7273 48546 7363
rect 45838 7213 45880 7273
rect 47877 7213 48546 7273
rect 45838 7160 48546 7213
rect 48816 7160 48855 8280
rect 45838 7127 48855 7160
rect 49073 -824 49433 16269
rect 45847 -888 49433 -824
rect 45847 -946 45884 -888
rect 48005 -946 49433 -888
rect 45847 -1007 49433 -946
rect 4254 -1161 19726 -1041
rect 49073 -1043 49433 -1007
rect 49553 26791 49913 35112
rect 49553 25616 49574 26791
rect 49888 25616 49913 26791
rect 49553 8284 49913 25616
rect 49553 7150 49576 8284
rect 49888 7150 49913 8284
rect 49553 -1043 49913 7150
<< via3 >>
rect 30 33050 220 34198
rect 1132 4936 1344 6296
<< metal4 >>
rect 1063 6296 1663 6318
rect 1063 4936 1132 6296
rect 1344 4936 1663 6296
rect 1063 4918 1663 4936
rect 1063 3031 1663 4716
rect 1063 1195 1663 2880
rect 1063 -564 1663 996
use bias_generator_fe  bias_generator_fe_0
timestamp 1720036258
transform 1 0 -35 0 1 -1186
box 1072 0 45976 8863
use bias_generator_idac_be  bias_generator_idac_be_0
timestamp 1720037216
transform 1 0 -89608 0 1 9596
box 88536 -10736 139522 25480
<< labels >>
flabel metal1 1037 3371 1437 3439 0 FreeSans 480 0 0 0 ena
port 53 nsew
flabel metal1 1037 4999 1437 5067 0 FreeSans 480 0 0 0 ref_sel_vbg
port 52 nsew
flabel metal1 435 7250 754 7371 0 FreeSans 640 0 0 0 vbg
port 54 nsew
flabel metal4 1063 -564 1547 996 0 FreeSans 3200 90 0 0 dvss
port 50 nsew
flabel metal4 1063 1195 1663 2880 0 FreeSans 3200 90 0 0 avss
port 12 nsew
flabel metal4 1063 3031 1663 4716 0 FreeSans 3200 90 0 0 avdd
port 59 nsew
flabel metal4 s 1063 4918 1663 6318 0 FreeSans 3200 90 0 0 dvdd
port 58 n
flabel metal3 49073 -1043 49433 -118 0 FreeSans 1600 90 0 0 snk_out
port 60 nsew
flabel metal3 49553 -1043 49913 -114 0 FreeSans 1600 90 0 0 src_out
port 61 nsew
flabel metal2 142 34487 182 34862 0 FreeSans 400 270 0 0 din[0]
port 22 nsew
flabel metal2 262 34487 302 34862 0 FreeSans 400 270 0 0 din[1]
port 23 nsew
flabel metal2 382 34487 422 34862 0 FreeSans 400 270 0 0 din[2]
port 21 nsew
flabel metal2 502 34487 542 34862 0 FreeSans 400 270 0 0 din[3]
port 20 nsew
flabel metal2 2734 34487 2774 34862 0 FreeSans 400 270 0 0 din[4]
port 25 nsew
flabel metal2 2854 34487 2894 34862 0 FreeSans 400 270 0 0 din[5]
port 24 nsew
flabel metal2 2970 34487 3010 34862 0 FreeSans 400 270 0 0 din[6]
port 16 nsew
flabel metal2 3094 34462 3134 34862 0 FreeSans 400 270 0 0 din[7]
port 26 nsew
flabel metal3 4254 -1161 4658 -1041 0 FreeSans 1120 0 0 0 ref_in
port 62 nsew
<< end >>
