magic
tech sky130A
magscale 1 2
timestamp 1717105881
<< error_s >>
rect 139295 4795 139298 4806
rect 139295 4778 139323 4795
rect 106922 4738 106931 4747
rect 106913 4729 106927 4738
rect 106922 4663 106927 4729
rect 106913 4654 106927 4663
rect 106922 4645 106931 4654
rect 106922 4379 106927 4463
rect 106776 925 107676 1825
rect 116972 278 117000 326
<< dnwell >>
rect 106776 719 138229 8571
<< nwell >>
rect 106776 8365 138338 8680
rect 138023 925 138338 8365
rect 106776 610 138338 925
<< pwell >>
rect 108895 925 108983 947
<< mvpsubdiff >>
rect 106842 8770 106922 8804
rect 138398 8770 138458 8804
rect 138424 8744 138458 8770
rect 139072 8182 139132 8216
rect 147424 8182 147484 8216
rect 139072 8156 139106 8182
rect 139072 1252 139106 1278
rect 147450 8156 147484 8182
rect 147450 1252 147484 1278
rect 139072 1218 139132 1252
rect 147424 1218 147484 1252
rect 138424 498 138458 524
rect 106842 464 106922 498
rect 138398 464 138458 498
<< mvnsubdiff >>
rect 106842 8594 138272 8614
rect 106842 8560 106922 8594
rect 138192 8560 138272 8594
rect 106842 8540 138272 8560
rect 138198 8534 138272 8540
rect 138198 756 138218 8534
rect 138252 756 138272 8534
rect 138198 750 138272 756
rect 106842 730 138272 750
rect 106842 696 106922 730
rect 138192 696 138272 730
rect 106842 676 138272 696
<< mvpsubdiffcont >>
rect 106922 8770 138398 8804
rect 138424 524 138458 8744
rect 139132 8182 147424 8216
rect 139072 1278 139106 8156
rect 147450 1278 147484 8156
rect 139132 1218 147424 1252
rect 106922 464 138398 498
<< mvnsubdiffcont >>
rect 106922 8560 138192 8594
rect 138218 756 138252 8534
rect 106922 696 138192 730
<< locali >>
rect 106842 8770 106922 8804
rect 138398 8770 138458 8804
rect 106842 8755 138458 8770
rect 106842 8671 138360 8755
rect 106850 8560 106922 8594
rect 138192 8560 138252 8594
rect 106850 8534 138252 8560
rect 106850 8529 138218 8534
rect 106850 8375 138128 8529
rect 138081 909 138128 8375
rect 106842 752 138128 909
rect 138187 756 138218 8529
rect 138187 752 138252 756
rect 106842 730 138252 752
rect 106842 696 106922 730
rect 138192 696 138252 730
rect 138316 610 138360 8671
rect 106842 523 138360 610
rect 106842 464 106922 523
rect 138307 514 138360 523
rect 138412 8744 138458 8755
rect 138412 524 138424 8744
rect 138458 8182 139132 8216
rect 147424 8182 147484 8216
rect 138458 8156 147484 8182
rect 138458 8019 139072 8156
rect 138458 1278 139072 1414
rect 139106 8094 147450 8156
rect 139106 1340 139189 8094
rect 139871 7594 139918 7660
rect 142463 7594 142510 7660
rect 145055 7594 145102 7660
rect 141509 6766 141679 6782
rect 141509 6664 141525 6766
rect 141658 6664 141679 6766
rect 141509 6648 141679 6664
rect 144101 6766 144271 6782
rect 144101 6664 144117 6766
rect 144250 6664 144271 6766
rect 144101 6648 144271 6664
rect 146693 6766 146863 6782
rect 146693 6664 146709 6766
rect 146842 6664 146863 6766
rect 146693 6648 146863 6664
rect 139871 5966 139918 6032
rect 142463 5966 142510 6032
rect 145055 5966 145102 6032
rect 141509 5138 141679 5154
rect 141509 5036 141525 5138
rect 141658 5036 141679 5138
rect 141509 5020 141679 5036
rect 144101 5138 144271 5154
rect 144101 5036 144117 5138
rect 144250 5036 144271 5138
rect 144101 5020 144271 5036
rect 146693 5138 146863 5154
rect 146693 5036 146709 5138
rect 146842 5036 146863 5138
rect 146693 5020 146863 5036
rect 142463 4338 142510 4404
rect 145055 4338 145102 4404
rect 141509 3510 141679 3526
rect 141509 3408 141525 3510
rect 141658 3408 141679 3510
rect 141509 3392 141679 3408
rect 144101 3510 144271 3526
rect 144101 3408 144117 3510
rect 144250 3408 144271 3510
rect 144101 3392 144271 3408
rect 146693 3510 146863 3526
rect 146693 3408 146709 3510
rect 146842 3408 146863 3510
rect 146693 3392 146863 3408
rect 142463 2710 142510 2776
rect 145055 2710 145102 2776
rect 141509 1882 141679 1898
rect 141509 1780 141525 1882
rect 141658 1780 141679 1882
rect 141509 1764 141679 1780
rect 144101 1882 144271 1898
rect 144101 1780 144117 1882
rect 144250 1780 144271 1882
rect 144101 1764 144271 1780
rect 146693 1882 146863 1898
rect 146693 1780 146709 1882
rect 146842 1780 146863 1882
rect 146693 1764 146863 1780
rect 147356 1340 147450 8094
rect 139106 1278 147450 1340
rect 138458 1252 147484 1278
rect 138458 1218 139132 1252
rect 147424 1218 147484 1252
rect 138458 1217 139161 1218
rect 138412 514 138458 524
rect 138307 498 138458 514
rect 138398 464 138458 498
<< viali >>
rect 138128 752 138187 8529
rect 106922 498 138307 523
rect 138360 514 138412 8755
rect 139537 7624 139583 7803
rect 142129 7624 142175 7803
rect 144721 7624 144767 7803
rect 141525 6664 141658 6766
rect 144117 6664 144250 6766
rect 146709 6664 146842 6766
rect 139537 5996 139583 6175
rect 142129 5996 142175 6175
rect 144721 5996 144767 6175
rect 141525 5036 141658 5138
rect 144117 5036 144250 5138
rect 146709 5036 146842 5138
rect 142129 4368 142175 4547
rect 144721 4368 144767 4547
rect 139918 4060 139966 4291
rect 141525 3408 141658 3510
rect 144117 3408 144250 3510
rect 146709 3408 146842 3510
rect 142129 2740 142175 2919
rect 144721 2740 144767 2919
rect 139918 2432 139966 2663
rect 141525 1780 141658 1882
rect 144117 1780 144250 1882
rect 146709 1780 146842 1882
rect 106922 479 138307 498
<< metal1 >>
rect 138332 8755 138448 8797
rect 138093 8529 138231 8580
rect 138093 6299 138128 8529
rect 138187 6299 138231 8529
rect 138093 4657 138108 6299
rect 138215 4657 138231 6299
rect 138093 752 138128 4657
rect 138187 752 138231 4657
rect 138093 705 138231 752
rect 138332 542 138360 8755
rect 138412 2512 138448 8755
rect 139334 8031 147268 8045
rect 139334 7872 140023 8031
rect 141298 7872 147268 8031
rect 139520 7815 139584 7816
rect 142116 7815 142180 7816
rect 139520 7814 139589 7815
rect 139520 7784 139526 7814
rect 139578 7803 139589 7814
rect 139480 7744 139526 7784
rect 139520 7614 139526 7744
rect 139583 7624 139589 7803
rect 139578 7614 139589 7624
rect 142116 7814 142181 7815
rect 142116 7614 142122 7814
rect 142174 7803 142181 7814
rect 142175 7624 142181 7803
rect 142174 7614 142181 7624
rect 139530 7612 139589 7614
rect 142122 7612 142181 7614
rect 144712 7814 144776 7816
rect 144712 7614 144718 7814
rect 144770 7614 144776 7814
rect 144712 7612 144776 7614
rect 142140 7529 142180 7612
rect 144728 7600 144768 7612
rect 139334 7066 142601 7239
rect 143880 7066 147257 7239
rect 139334 6946 145336 7003
rect 141509 6766 141679 6782
rect 141509 6664 141525 6766
rect 141658 6664 141679 6766
rect 141509 6648 141679 6664
rect 144101 6766 144271 6782
rect 144101 6664 144117 6766
rect 144250 6664 144271 6766
rect 144101 6648 144271 6664
rect 146693 6766 146863 6782
rect 146693 6664 146709 6766
rect 146842 6664 146863 6766
rect 146693 6648 146863 6664
rect 139334 6249 140026 6422
rect 141296 6249 147257 6422
rect 139520 6187 139584 6188
rect 139520 6186 139589 6187
rect 139520 6156 139526 6186
rect 139578 6175 139589 6186
rect 139490 6116 139526 6156
rect 139520 5986 139526 6116
rect 139583 5996 139589 6175
rect 139578 5986 139589 5996
rect 142116 6186 142182 6188
rect 144714 6186 144773 6187
rect 142116 5986 142122 6186
rect 142174 6175 142182 6186
rect 142175 5996 142182 6175
rect 142174 5986 142182 5996
rect 144712 5986 144718 6186
rect 144770 5986 144776 6186
rect 139530 5984 139589 5986
rect 142122 5984 142181 5986
rect 144712 5984 144776 5986
rect 142140 5901 142180 5984
rect 144728 5980 144768 5984
rect 139334 5438 142597 5611
rect 143876 5438 147274 5611
rect 139334 5318 145336 5375
rect 141509 5138 141679 5154
rect 141509 5036 141525 5138
rect 141658 5036 141679 5138
rect 141509 5020 141679 5036
rect 144101 5138 144271 5154
rect 144101 5036 144117 5138
rect 144250 5036 144271 5138
rect 144101 5020 144271 5036
rect 146693 5138 146863 5154
rect 146693 5036 146709 5138
rect 146842 5036 146863 5138
rect 146693 5020 146863 5036
rect 139295 4778 139298 4795
rect 139334 4622 140024 4795
rect 141294 4622 147246 4795
rect 142116 4559 142180 4560
rect 142116 4558 142181 4559
rect 144714 4558 144773 4559
rect 142116 4528 142122 4558
rect 142174 4547 142181 4558
rect 138822 4168 138828 4368
rect 138880 4328 139967 4368
rect 142116 4358 142122 4488
rect 142175 4368 142181 4547
rect 142174 4358 142181 4368
rect 142122 4356 142181 4358
rect 144712 4358 144718 4558
rect 144770 4358 144776 4558
rect 144712 4356 144776 4358
rect 144728 4350 144768 4356
rect 138880 4168 138886 4328
rect 139927 4297 139967 4328
rect 139906 4291 139982 4297
rect 139906 4060 139918 4291
rect 139966 4060 139982 4291
rect 139906 4054 139982 4060
rect 139334 3822 142601 3995
rect 143880 3822 147263 3995
rect 139334 3690 145336 3747
rect 141509 3510 141679 3526
rect 141509 3408 141525 3510
rect 141658 3408 141679 3510
rect 141509 3392 141679 3408
rect 144101 3510 144271 3526
rect 144101 3408 144117 3510
rect 144250 3408 144271 3510
rect 144101 3392 144271 3408
rect 146693 3510 146863 3526
rect 146693 3408 146709 3510
rect 146842 3408 146863 3510
rect 146693 3392 146863 3408
rect 139334 3000 140028 3173
rect 141298 3000 147230 3173
rect 142116 2930 142182 2932
rect 144714 2930 144773 2931
rect 142116 2900 142122 2930
rect 142174 2919 142182 2930
rect 138932 2540 138938 2740
rect 138990 2700 139963 2740
rect 142116 2730 142122 2860
rect 142175 2740 142182 2919
rect 142174 2730 142182 2740
rect 144712 2730 144718 2930
rect 144770 2730 144776 2930
rect 142122 2728 142181 2730
rect 144712 2728 144776 2730
rect 144728 2710 144768 2728
rect 138990 2540 138996 2700
rect 139923 2669 139963 2700
rect 139906 2663 139979 2669
rect 138412 2481 138622 2512
rect 138593 1342 138622 2481
rect 139906 2432 139918 2663
rect 139966 2432 139979 2663
rect 139906 2426 139979 2432
rect 139334 2183 142601 2356
rect 143880 2183 147274 2356
rect 139334 2062 145336 2119
rect 141509 1882 141679 1898
rect 141509 1780 141525 1882
rect 141658 1780 141679 1882
rect 141509 1764 141679 1780
rect 144101 1882 144271 1898
rect 144101 1780 144117 1882
rect 144250 1780 144271 1882
rect 144101 1764 144271 1780
rect 146693 1882 146863 1898
rect 146693 1780 146709 1882
rect 146842 1780 146863 1882
rect 146693 1764 146863 1780
rect 139334 1461 140021 1539
rect 141293 1461 147196 1539
rect 106842 523 138360 542
rect 106842 479 106922 523
rect 138307 514 138360 523
rect 138412 1310 138622 1342
rect 138412 514 138448 1310
rect 138307 479 138448 514
rect 106842 464 138448 479
<< via1 >>
rect 138108 4657 138128 6299
rect 138128 4657 138187 6299
rect 138187 4657 138215 6299
rect 140023 7868 141298 8031
rect 139526 7803 139578 7814
rect 139526 7624 139537 7803
rect 139537 7624 139578 7803
rect 139526 7614 139578 7624
rect 142122 7803 142174 7814
rect 142122 7624 142129 7803
rect 142129 7624 142174 7803
rect 142122 7614 142174 7624
rect 144718 7803 144770 7814
rect 144718 7624 144721 7803
rect 144721 7624 144767 7803
rect 144767 7624 144770 7803
rect 144718 7614 144770 7624
rect 142601 7047 143880 7264
rect 145336 6946 146330 7003
rect 141525 6664 141658 6766
rect 144117 6664 144250 6766
rect 146709 6664 146842 6766
rect 140026 6229 141296 6444
rect 139526 6175 139578 6186
rect 139526 5996 139537 6175
rect 139537 5996 139578 6175
rect 139526 5986 139578 5996
rect 142122 6175 142174 6186
rect 142122 5996 142129 6175
rect 142129 5996 142174 6175
rect 142122 5986 142174 5996
rect 144718 6175 144770 6186
rect 144718 5996 144721 6175
rect 144721 5996 144767 6175
rect 144767 5996 144770 6175
rect 144718 5986 144770 5996
rect 142597 5420 143876 5637
rect 145336 5318 146330 5375
rect 141525 5036 141658 5138
rect 144117 5036 144250 5138
rect 146709 5036 146842 5138
rect 140024 4609 141294 4824
rect 142122 4547 142174 4558
rect 138828 4168 138880 4368
rect 142122 4368 142129 4547
rect 142129 4368 142174 4547
rect 142122 4358 142174 4368
rect 144718 4547 144770 4558
rect 144718 4368 144721 4547
rect 144721 4368 144767 4547
rect 144767 4368 144770 4547
rect 144718 4358 144770 4368
rect 142601 3789 143880 4006
rect 145336 3690 146330 3747
rect 141525 3408 141658 3510
rect 144117 3408 144250 3510
rect 146709 3408 146842 3510
rect 140028 2976 141298 3191
rect 142122 2919 142174 2930
rect 138938 2540 138990 2740
rect 142122 2740 142129 2919
rect 142129 2740 142174 2919
rect 142122 2730 142174 2740
rect 144718 2919 144770 2930
rect 144718 2740 144721 2919
rect 144721 2740 144767 2919
rect 144767 2740 144770 2919
rect 144718 2730 144770 2740
rect 138379 1342 138412 2481
rect 138412 1342 138593 2481
rect 142601 2163 143880 2380
rect 145336 2062 146330 2119
rect 141525 1780 141658 1882
rect 144117 1780 144250 1882
rect 146709 1780 146842 1882
rect 140021 1448 141293 1563
<< metal2 >>
rect 127394 9730 145084 9778
rect 127394 9346 127442 9730
rect 117318 9298 127442 9346
rect 127550 9634 144898 9682
rect 117318 9138 117366 9298
rect 127550 9254 127598 9634
rect 106922 9090 117366 9138
rect 117506 9206 127598 9254
rect 127696 9538 144764 9586
rect 107110 8735 112834 8967
rect 113161 8735 117368 8967
rect 117506 8660 117554 9206
rect 127696 9134 127744 9538
rect 123920 9086 127744 9134
rect 128202 9442 144628 9490
rect 117754 8735 121402 8967
rect 121729 8735 123820 8967
rect 123920 8660 123968 9086
rect 124170 8735 126662 8967
rect 126989 8735 128064 8967
rect 128202 8660 128250 9442
rect 130336 9346 142486 9394
rect 128539 8735 129832 8967
rect 130159 8735 130186 8967
rect 130336 8660 130384 9346
rect 134516 9250 142330 9298
rect 134516 9114 134564 9250
rect 132658 9066 134564 9114
rect 134708 9154 142168 9202
rect 130685 8735 131924 8967
rect 132251 8735 132590 8967
rect 132658 8660 132706 9066
rect 132825 8735 134016 8967
rect 134343 8735 134640 8967
rect 134708 8660 134756 9154
rect 107270 8428 111939 8660
rect 112124 8428 117562 8660
rect 117926 8428 120507 8660
rect 120692 8428 123968 8660
rect 124197 8428 125767 8660
rect 125952 8428 128250 8660
rect 128617 8428 128937 8660
rect 129122 8428 130384 8660
rect 130721 8428 131029 8660
rect 131214 8612 132706 8660
rect 131214 8428 132590 8612
rect 132825 8428 133121 8660
rect 133306 8612 134756 8660
rect 134812 9058 142020 9106
rect 134812 8658 134860 9058
rect 134929 8735 135568 8967
rect 135895 8735 135909 8967
rect 135981 8735 135997 8967
rect 136169 8735 136203 8967
rect 136506 8735 136678 8967
rect 136895 8735 137113 8967
rect 134929 8658 135213 8660
rect 133306 8428 134640 8612
rect 134812 8610 135213 8658
rect 134929 8428 135213 8610
rect 135398 8428 135858 8660
rect 135981 8428 136339 8660
rect 136524 8428 136549 8660
rect 136693 8428 137022 8660
rect 137197 8520 137292 8660
rect 137197 8480 139572 8520
rect 137197 8428 137292 8480
rect 136494 8372 136534 8428
rect 139362 8372 139402 8376
rect 136494 8332 139402 8372
rect 106866 8027 137616 8265
rect 106866 7696 106988 7930
rect 137608 7696 137655 7930
rect 137910 7696 137939 7930
rect 139362 7384 139402 8332
rect 139532 7824 139572 8480
rect 140008 8031 141311 8086
rect 140008 7868 140023 8031
rect 141298 7868 141311 8031
rect 139526 7814 139578 7824
rect 139526 7606 139578 7614
rect 139362 7344 139572 7384
rect 106866 6696 137616 6930
rect 106866 6695 106986 6696
rect 138079 6299 138270 6322
rect 106922 5692 137616 5926
rect 137608 4638 137654 4872
rect 137909 4638 137938 4872
rect 138079 4657 138108 6299
rect 138215 4657 138270 6299
rect 139532 6196 139572 7344
rect 140008 6444 141311 7868
rect 141980 7194 142020 9058
rect 142128 7824 142168 9154
rect 142122 7814 142174 7824
rect 142122 7606 142174 7614
rect 141980 7154 142168 7194
rect 141509 6766 141679 6782
rect 141509 6664 141525 6766
rect 141658 6739 141679 6766
rect 141658 6699 142039 6739
rect 141658 6664 141679 6699
rect 141509 6648 141679 6664
rect 140008 6229 140026 6444
rect 141296 6229 141311 6444
rect 139526 6186 139578 6196
rect 139526 5978 139578 5986
rect 138079 4638 138270 4657
rect 140008 4824 141311 6229
rect 141509 5138 141679 5154
rect 141509 5036 141525 5138
rect 141658 5097 141679 5138
rect 141658 5057 141919 5097
rect 141658 5036 141679 5057
rect 141509 5020 141679 5036
rect 140008 4609 140024 4824
rect 141294 4609 141311 4824
rect 106866 4463 108079 4480
rect 106866 4379 106922 4463
rect 106866 4377 107192 4379
rect 106866 4242 108079 4377
rect 138828 4368 138880 4376
rect 138828 4162 138880 4168
rect 106922 3218 137597 3456
rect 138358 2481 138622 2512
rect 106922 2234 137589 2472
rect 106866 1246 137597 1484
rect 138358 1342 138379 2481
rect 138593 1342 138622 2481
rect 138358 1310 138622 1342
rect 138834 1172 138874 4162
rect 140008 3191 141311 4609
rect 141509 3510 141679 3526
rect 141509 3408 141525 3510
rect 141658 3474 141679 3510
rect 141658 3434 141803 3474
rect 141658 3408 141679 3434
rect 141509 3392 141679 3408
rect 140008 2976 140028 3191
rect 141298 2976 141311 3191
rect 138938 2740 138990 2748
rect 138938 2534 138990 2540
rect 136210 1132 138874 1172
rect 136210 1037 136250 1132
rect 106866 849 120004 1037
rect 120189 849 136250 1037
rect 136690 849 137068 1037
rect 137185 972 137300 1037
rect 138944 972 138984 2534
rect 140008 2485 141311 2976
rect 140008 1563 140035 2485
rect 141277 1563 141311 2485
rect 141509 1882 141679 1898
rect 141509 1780 141525 1882
rect 141658 1780 141679 1882
rect 141509 1764 141679 1780
rect 140008 1448 140021 1563
rect 141293 1448 141311 1563
rect 140008 1340 140035 1448
rect 141277 1340 141311 1448
rect 140008 1300 141311 1340
rect 137185 932 138984 972
rect 137185 849 137300 932
rect 106866 593 120899 781
rect 121226 593 136081 781
rect 136525 593 136680 781
rect 136862 593 137135 781
rect 141639 678 141679 1764
rect 141759 1096 141803 3434
rect 141763 678 141803 1096
rect 141879 678 141919 5057
rect 141999 678 142039 6699
rect 142128 6196 142168 7154
rect 142122 6186 142174 6196
rect 142122 5978 142174 5986
rect 142290 5302 142330 9250
rect 142128 5262 142330 5302
rect 142128 4568 142168 5262
rect 142122 4558 142174 4568
rect 142122 4350 142174 4358
rect 142446 4076 142486 9346
rect 142128 4036 142486 4076
rect 142588 7264 143893 8101
rect 142588 7047 142601 7264
rect 143880 7047 143893 7264
rect 144588 7178 144628 9442
rect 144724 7824 144764 9538
rect 144718 7814 144770 7824
rect 144718 7606 144770 7614
rect 144588 7138 144764 7178
rect 142588 6280 143893 7047
rect 144101 6766 144271 6782
rect 144101 6664 144117 6766
rect 144250 6739 144271 6766
rect 144250 6699 144631 6739
rect 144250 6664 144271 6699
rect 144101 6648 144271 6664
rect 142588 5637 142647 6280
rect 143849 5637 143893 6280
rect 142588 5420 142597 5637
rect 143876 5420 143893 5637
rect 142588 4689 142647 5420
rect 143849 4689 143893 5420
rect 144101 5138 144271 5154
rect 144101 5036 144117 5138
rect 144250 5097 144271 5138
rect 144250 5057 144511 5097
rect 144250 5036 144271 5057
rect 144101 5020 144271 5036
rect 142128 2940 142168 4036
rect 142588 4006 143893 4689
rect 142588 3789 142601 4006
rect 143880 3789 143893 4006
rect 142122 2930 142174 2940
rect 142122 2722 142174 2730
rect 142588 2380 143893 3789
rect 144101 3510 144271 3526
rect 144101 3408 144117 3510
rect 144250 3474 144271 3510
rect 144250 3434 144391 3474
rect 144250 3408 144271 3434
rect 144101 3392 144271 3408
rect 142588 2163 142601 2380
rect 143880 2163 143893 2380
rect 142588 1390 143893 2163
rect 144101 1882 144271 1898
rect 144101 1780 144117 1882
rect 144250 1780 144271 1882
rect 144101 1764 144271 1780
rect 144231 678 144271 1764
rect 144351 678 144391 3434
rect 144471 678 144511 5057
rect 144591 678 144631 6699
rect 144724 6196 144764 7138
rect 144718 6186 144770 6196
rect 144718 5978 144770 5986
rect 144858 5870 144898 9634
rect 144724 5830 144898 5870
rect 144724 4568 144764 5830
rect 144718 4558 144770 4568
rect 144718 4350 144770 4358
rect 145044 4090 145084 9730
rect 144724 4050 145084 4090
rect 145336 7851 146330 8094
rect 145336 7003 145367 7851
rect 146299 7003 146330 7851
rect 145336 6713 145367 6946
rect 146299 6713 146330 6946
rect 145336 5375 146330 6713
rect 146693 6766 146863 6782
rect 146693 6664 146709 6766
rect 146842 6739 146863 6766
rect 146842 6699 147223 6739
rect 146842 6664 146863 6699
rect 146693 6648 146863 6664
rect 144724 2940 144764 4050
rect 145336 3747 146330 5318
rect 146693 5138 146863 5154
rect 146693 5036 146709 5138
rect 146842 5097 146863 5138
rect 146842 5057 147103 5097
rect 146842 5036 146863 5057
rect 146693 5020 146863 5036
rect 144718 2930 144770 2940
rect 144718 2722 144770 2730
rect 145336 2119 146330 3690
rect 146693 3510 146863 3526
rect 146693 3408 146709 3510
rect 146842 3474 146863 3510
rect 146842 3434 146983 3474
rect 146842 3408 146863 3434
rect 146693 3392 146863 3408
rect 145336 1301 146330 2062
rect 146693 1882 146863 1898
rect 146693 1780 146709 1882
rect 146842 1780 146863 1882
rect 146693 1764 146863 1780
rect 146823 1146 146863 1764
rect 146943 678 146983 3434
rect 147063 678 147103 5057
rect 147183 678 147223 6699
rect 116972 278 116978 326
<< via2 >>
rect 112834 8735 113161 8967
rect 121402 8735 121729 8967
rect 126662 8735 126989 8967
rect 129832 8735 130159 8967
rect 131924 8735 132251 8967
rect 134016 8735 134343 8967
rect 111939 8428 112124 8660
rect 120507 8428 120692 8660
rect 125767 8428 125952 8660
rect 128937 8428 129122 8660
rect 131029 8428 131214 8660
rect 133121 8428 133306 8660
rect 135568 8735 135895 8967
rect 135997 8735 136169 8967
rect 136678 8735 136895 8967
rect 135213 8428 135398 8660
rect 136339 8428 136524 8660
rect 137022 8428 137197 8660
rect 137655 7696 137910 7930
rect 106922 4654 137146 4738
rect 137654 4638 137909 4872
rect 138108 4657 138215 6299
rect 106922 4379 137147 4463
rect 107192 4377 109062 4379
rect 138379 1342 138593 2481
rect 120004 849 120189 1037
rect 137068 849 137185 1037
rect 140035 1563 141277 2485
rect 140035 1448 141277 1563
rect 140035 1340 141277 1448
rect 120899 593 121226 781
rect 136680 593 136862 781
rect 142647 5637 143849 6280
rect 142647 5420 143849 5637
rect 142647 4689 143849 5420
rect 145367 7003 146299 7851
rect 145367 6946 146299 7003
rect 145367 6713 146299 6946
<< metal3 >>
rect 111922 8660 112143 9465
rect 112817 8967 113179 9465
rect 112817 8735 112834 8967
rect 113161 8735 113179 8967
rect 112817 8714 113179 8735
rect 111922 8428 111939 8660
rect 112124 8428 112143 8660
rect 111922 8390 112143 8428
rect 120490 8660 120711 9466
rect 121385 8967 121747 9465
rect 121385 8735 121402 8967
rect 121729 8735 121747 8967
rect 121385 8714 121747 8735
rect 120490 8428 120507 8660
rect 120692 8428 120711 8660
rect 120490 8390 120711 8428
rect 125750 8660 125971 9465
rect 126645 8967 127003 9465
rect 126645 8735 126662 8967
rect 126989 8735 127003 8967
rect 126645 8714 127003 8735
rect 125750 8428 125767 8660
rect 125952 8428 125971 8660
rect 125750 8390 125971 8428
rect 128920 8660 129141 9465
rect 129815 8967 130173 9465
rect 129815 8735 129832 8967
rect 130159 8735 130173 8967
rect 129815 8714 130173 8735
rect 128920 8428 128937 8660
rect 129122 8428 129141 8660
rect 128920 8390 129141 8428
rect 131012 8660 131233 9465
rect 131907 8967 132265 9465
rect 131907 8735 131924 8967
rect 132251 8735 132265 8967
rect 131907 8714 132265 8735
rect 131012 8428 131029 8660
rect 131214 8428 131233 8660
rect 131012 8390 131233 8428
rect 133104 8660 133325 9465
rect 133999 8967 134357 9465
rect 133999 8735 134016 8967
rect 134343 8735 134357 8967
rect 133999 8714 134357 8735
rect 133104 8428 133121 8660
rect 133306 8428 133325 8660
rect 133104 8390 133325 8428
rect 135196 8660 135417 9465
rect 135551 8967 135909 9465
rect 135551 8735 135568 8967
rect 135895 8735 135909 8967
rect 135551 8714 135909 8735
rect 135980 8967 136219 9465
rect 135980 8735 135997 8967
rect 136169 8735 136219 8967
rect 135980 8714 136219 8735
rect 135196 8428 135213 8660
rect 135398 8428 135417 8660
rect 135196 8390 135417 8428
rect 136322 8660 136543 9465
rect 136664 8967 136907 9466
rect 136664 8735 136678 8967
rect 136895 8735 136907 8967
rect 136664 8715 136907 8735
rect 136322 8428 136339 8660
rect 136524 8428 136543 8660
rect 136322 8390 136543 8428
rect 137011 8660 137210 9467
rect 137011 8428 137022 8660
rect 137197 8428 137210 8660
rect 137011 8408 137210 8428
rect 137642 7930 137920 7967
rect 137642 7696 137655 7930
rect 137910 7696 137920 7930
rect 137642 4872 137920 7696
rect 145336 7851 146329 7886
rect 145336 6713 145367 7851
rect 146299 6713 146329 7851
rect 145336 6684 146329 6713
rect 106922 4827 137654 4872
rect 137147 4653 137654 4827
rect 106922 4638 137654 4653
rect 137909 4638 137920 4872
rect 138079 6299 138248 6321
rect 138079 4657 138108 6299
rect 138215 4657 138248 6299
rect 138079 4638 138248 4657
rect 142588 6280 143894 6323
rect 142588 4689 142647 6280
rect 143849 4689 143894 6280
rect 106922 4464 137539 4480
rect 137147 4290 137539 4464
rect 106922 4288 107192 4290
rect 109062 4288 137539 4290
rect 106922 4242 137539 4288
rect 137642 1254 137920 4638
rect 142588 4636 143894 4689
rect 138358 2481 138622 2512
rect 138358 1342 138379 2481
rect 138593 1342 138622 2481
rect 138358 1310 138622 1342
rect 140009 2485 141309 2513
rect 140009 1340 140035 2485
rect 141277 1340 141309 2485
rect 140009 1313 141309 1340
rect 119987 1037 120208 1076
rect 119987 849 120004 1037
rect 120189 849 120208 1037
rect 119987 1 120208 849
rect 137060 1037 137194 1053
rect 137060 849 137068 1037
rect 137185 849 137194 1037
rect 120882 781 121244 803
rect 120882 593 120899 781
rect 121226 593 121244 781
rect 120882 1 121244 593
rect 136670 781 136875 800
rect 136670 593 136680 781
rect 136862 593 136875 781
rect 136670 193 136875 593
rect 137060 195 137194 849
<< via3 >>
rect 145367 6713 146299 7851
rect 106922 4738 137147 4827
rect 106922 4654 137146 4738
rect 137146 4654 137147 4738
rect 106922 4653 137147 4654
rect 138108 4657 138215 6299
rect 142647 4689 143849 6280
rect 106922 4463 137147 4464
rect 106922 4379 137147 4463
rect 106922 4377 107192 4379
rect 107192 4377 109062 4379
rect 109062 4377 137147 4379
rect 106922 4290 137147 4377
rect 107192 4288 109062 4290
rect 138379 1342 138593 2481
rect 140035 1340 141277 2485
<< metal4 >>
rect 138356 7851 147485 7883
rect 138356 6713 145367 7851
rect 146299 6713 147485 7851
rect 138356 6683 147485 6713
rect 106865 6299 147485 6320
rect 106865 4827 138108 6299
rect 106865 4653 106922 4827
rect 137147 4657 138108 4827
rect 138215 6280 147485 6299
rect 138215 4689 142647 6280
rect 143849 4689 147485 6280
rect 138215 4657 147485 4689
rect 137147 4653 147485 4657
rect 106865 4635 147485 4653
rect 106866 4464 147485 4484
rect 106866 4290 106922 4464
rect 137147 4290 147485 4464
rect 106866 4288 107192 4290
rect 109062 4288 147485 4290
rect 106866 2799 147485 4288
rect 138356 2485 147485 2511
rect 138356 2481 140035 2485
rect 138356 1342 138379 2481
rect 138593 1342 140035 2481
rect 138356 1340 140035 1342
rect 141277 1340 147485 2485
rect 138356 1311 147485 1340
use bias_nstack  bias_nstack_0
array 0 56 -534 0 0 -3895
timestamp 1717035242
transform -1 0 110949 0 -1 1620
box 3258 -2860 3926 1035
use bias_pstack  bias_pstack_0
array 0 56 534 0 0 -4355
timestamp 1717035242
transform 1 0 104996 0 -1 5026
box 1986 -3967 2714 388
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_3 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform -1 0 145080 0 1 1458
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_5
timestamp 1715205430
transform -1 0 145080 0 1 6342
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_6
timestamp 1715205430
transform -1 0 145080 0 1 4714
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_7
timestamp 1715205430
transform -1 0 145080 0 1 3086
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_8
timestamp 1715205430
transform -1 0 142488 0 1 1458
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_9
timestamp 1715205430
transform -1 0 142488 0 1 4714
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_10
timestamp 1715205430
transform -1 0 142488 0 1 3086
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_11
timestamp 1715205430
transform -1 0 139896 0 1 1458
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_12
timestamp 1715205430
transform -1 0 142488 0 1 6342
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_13
timestamp 1715205430
transform -1 0 139896 0 1 6342
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_14
timestamp 1715205430
transform -1 0 139896 0 -1 3086
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_16
timestamp 1715205430
transform -1 0 139896 0 1 4714
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_17
timestamp 1715205430
transform -1 0 139896 0 1 3086
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_18
timestamp 1715205430
transform -1 0 139896 0 -1 4714
box -66 -43 450 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform -1 0 147288 0 -1 6342
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_1
timestamp 1715205430
transform -1 0 147288 0 -1 3086
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_2
timestamp 1715205430
transform -1 0 147288 0 -1 4714
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_3
timestamp 1715205430
transform -1 0 144696 0 1 1458
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_4
timestamp 1715205430
transform -1 0 147288 0 -1 7970
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_5
timestamp 1715205430
transform -1 0 144696 0 1 6342
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_6
timestamp 1715205430
transform -1 0 144696 0 1 4714
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_7
timestamp 1715205430
transform -1 0 144696 0 1 3086
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_8
timestamp 1715205430
transform -1 0 142104 0 1 1458
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_9
timestamp 1715205430
transform -1 0 142104 0 1 4714
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_10
timestamp 1715205430
transform -1 0 142104 0 1 3086
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_11
timestamp 1715205430
transform -1 0 139512 0 1 1458
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_12
timestamp 1715205430
transform -1 0 142104 0 1 6342
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_13
timestamp 1715205430
transform -1 0 139512 0 1 6342
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_14
timestamp 1715205430
transform -1 0 139512 0 -1 3086
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_16
timestamp 1715205430
transform -1 0 139512 0 1 4714
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_17
timestamp 1715205430
transform -1 0 139512 0 1 3086
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_18
timestamp 1715205430
transform -1 0 139512 0 -1 4714
box -66 -43 162 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform -1 0 145080 0 -1 3086
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_1
timestamp 1715205430
transform -1 0 139896 0 -1 7970
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_5
timestamp 1715205430
transform -1 0 145080 0 -1 7970
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_6
timestamp 1715205430
transform -1 0 145080 0 -1 6342
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_7
timestamp 1715205430
transform -1 0 145080 0 -1 4714
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_8
timestamp 1715205430
transform -1 0 142488 0 -1 4714
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_9
timestamp 1715205430
transform -1 0 142488 0 -1 3086
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_10
timestamp 1715205430
transform -1 0 142488 0 -1 7970
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_11
timestamp 1715205430
transform -1 0 142488 0 -1 6342
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_12
timestamp 1715205430
transform -1 0 139896 0 -1 6342
box -66 -43 546 897
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
array 0 2 -2592 0 3 1628
timestamp 1715205430
transform -1 0 142008 0 1 1458
box -66 -43 2178 1671
<< labels >>
flabel metal4 146885 6683 147485 7883 0 FreeSans 3200 90 0 0 dvdd
port 3 nsew
flabel metal4 146885 4635 147485 6320 0 FreeSans 3200 90 0 0 avdd
port 1 nsew
flabel metal4 146885 2799 147485 4484 0 FreeSans 3200 90 0 0 avss
port 2 nsew
flabel metal4 146885 1311 147485 2511 0 FreeSans 3200 90 0 0 dvss
port 4 nsew
flabel metal4 106866 2799 107099 4484 0 FreeSans 1600 90 0 0 avss
port 2 nsew
flabel metal4 106865 4635 107098 6320 0 FreeSans 1600 90 0 0 avdd
port 1 nsew
flabel metal3 136670 193 136875 335 0 FreeSans 1600 90 0 0 snk_test1
port 5 nsew
flabel metal3 136664 9225 136907 9466 0 FreeSans 1600 90 0 0 src_test1
port 6 nsew
flabel metal3 135980 9225 136219 9465 0 FreeSans 1600 90 0 0 src_50
port 7 nsew
flabel metal3 135551 9225 135909 9465 0 FreeSans 1600 90 0 0 src_100
port 8 nsew
flabel metal3 133999 9225 134357 9465 0 FreeSans 1600 90 0 0 src_200_2
port 9 nsew
flabel metal3 131907 9225 132265 9465 0 FreeSans 1600 90 0 0 src_200_1
port 10 nsew
flabel metal3 129815 9225 130173 9465 0 FreeSans 1600 90 0 0 src_200_0
port 11 nsew
flabel metal3 126645 9225 127003 9465 0 FreeSans 1600 90 0 0 src_400
port 12 nsew
flabel metal3 121385 9224 121747 9465 0 FreeSans 1600 90 0 0 src_600
port 13 nsew
flabel metal3 137060 195 137194 337 0 FreeSans 1600 90 0 0 ena_test1_3v3
flabel metal3 137011 9226 137210 9467 0 FreeSans 1600 90 0 0 enb_test1_3v3
flabel metal3 136322 9225 136543 9465 0 FreeSans 1600 90 0 0 enb_50_3v3
flabel metal3 135196 9225 135417 9465 0 FreeSans 1600 90 0 0 enb_100_3v3
flabel metal3 133104 9225 133325 9465 0 FreeSans 1600 90 0 0 enb_200_2_3v3
flabel metal3 131012 9225 131233 9465 0 FreeSans 1600 90 0 0 enb_200_1_3v3
flabel metal3 128920 9225 129141 9465 0 FreeSans 1600 90 0 0 enb_200_0_3v3
flabel metal3 125750 9225 125971 9465 0 FreeSans 1600 90 0 0 enb_400_3v3
flabel metal3 120490 9225 120711 9466 0 FreeSans 1600 90 0 0 enb_600_3v3
flabel metal3 119987 1 120208 189 0 FreeSans 1600 90 0 0 ena_test2_3v3
flabel metal3 111922 9224 112143 9465 0 FreeSans 1600 90 0 0 enb_1000_3v3
flabel metal3 112817 9224 113179 9465 0 FreeSans 1600 90 0 0 src_1000
port 14 nsew
flabel metal3 120882 1 121244 189 0 FreeSans 1600 90 0 0 snk_test2
port 15 nsew
flabel metal2 141763 678 141803 1053 0 FreeSans 400 90 0 0 ena_snk_test2
port 16 nsew
flabel metal3 146943 678 146983 1053 0 FreeSans 400 90 0 0 ena_src_1000
port 17 nsew
flabel metal3 147183 678 147223 1053 0 FreeSans 400 90 0 0 ena_src_600
port 18 nsew
flabel metal3 147063 678 147103 1053 0 FreeSans 400 90 0 0 ena_src_400
port 19 nsew
flabel metal3 144231 678 144271 1053 0 FreeSans 400 90 0 0 ena_src_200_0
port 20 nsew
flabel metal3 144351 678 144391 1053 0 FreeSans 400 90 0 0 ena_src_200_1
port 21 nsew
flabel metal3 144591 678 144631 1053 0 FreeSans 400 90 0 0 ena_src_200_2
port 22 nsew
flabel metal3 144471 678 144511 1053 0 FreeSans 400 90 0 0 ena_src_100
port 23 nsew
flabel metal3 141879 678 141919 1053 0 FreeSans 400 90 0 0 ena_src_50
port 24 nsew
flabel metal3 141999 678 142039 1053 0 FreeSans 400 90 0 0 ena_src_test1
port 25 nsew
flabel metal2 141639 678 141679 1078 0 FreeSans 400 90 0 0 ena_snk_test1
port 26 nsew
<< end >>
