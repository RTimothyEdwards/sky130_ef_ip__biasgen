magic
tech sky130A
magscale 1 2
timestamp 1747752274
<< error_s >>
rect 82746 925 83646 1825
<< dnwell >>
rect 82746 719 138229 8571
<< nwell >>
rect 82746 8365 138338 8680
rect 138023 925 138338 8365
rect 82746 610 138338 925
<< pwell >>
rect 108895 925 108983 947
<< mvpsubdiff >>
rect 82812 8770 83084 8804
rect 138398 8770 138458 8804
rect 138424 8744 138458 8770
rect 139072 8190 139132 8216
rect 139067 8182 139132 8190
rect 157792 8182 157852 8216
rect 139067 8156 157852 8182
rect 139067 1278 139072 8156
rect 139106 8098 157818 8156
rect 139106 7987 139175 8098
rect 157725 7987 157818 8098
rect 139106 7953 139429 7987
rect 157549 7953 157818 7987
rect 139106 6359 139175 7953
rect 157725 6359 157818 7953
rect 139106 6325 139429 6359
rect 157549 6325 157818 6359
rect 139106 4731 139175 6325
rect 157725 4731 157818 6325
rect 139106 4697 139429 4731
rect 157549 4697 157818 4731
rect 139106 3103 139175 4697
rect 157725 3103 157818 4697
rect 139106 3069 139429 3103
rect 157549 3069 157818 3103
rect 139106 1475 139175 3069
rect 157725 1475 157818 3069
rect 139106 1441 139429 1475
rect 157549 1441 157818 1475
rect 139106 1322 139175 1441
rect 157725 1322 157818 1441
rect 139106 1278 157818 1322
rect 139067 1252 157852 1278
rect 139067 1228 139132 1252
rect 139072 1218 139132 1228
rect 157792 1218 157852 1252
rect 138424 498 138458 524
rect 82812 464 83084 498
rect 138398 464 138458 498
<< mvnsubdiff >>
rect 82812 8594 138272 8614
rect 82812 8560 83084 8594
rect 138192 8560 138272 8594
rect 82812 8540 138272 8560
rect 138198 8534 138272 8540
rect 138198 756 138218 8534
rect 138252 756 138272 8534
rect 138198 750 138272 756
rect 82812 730 138272 750
rect 82812 696 83084 730
rect 138192 696 138272 730
rect 82812 676 138272 696
<< mvpsubdiffcont >>
rect 83084 8770 138398 8804
rect 138424 524 138458 8744
rect 139132 8182 157792 8216
rect 139072 1278 139106 8156
rect 157818 1278 157852 8156
rect 139132 1218 157792 1252
rect 83084 464 138398 498
<< mvnsubdiffcont >>
rect 83084 8560 138192 8594
rect 138218 756 138252 8534
rect 83084 696 138192 730
<< locali >>
rect 82812 8770 83084 8804
rect 138398 8770 138458 8804
rect 82812 8755 138458 8770
rect 82812 8671 138360 8755
rect 82820 8560 83084 8594
rect 138192 8560 138252 8594
rect 82820 8534 138252 8560
rect 82820 8529 138218 8534
rect 82820 8492 138128 8529
rect 82820 8426 137381 8492
rect 137531 8426 138128 8492
rect 82820 8375 138128 8426
rect 138081 909 138128 8375
rect 82812 752 138128 909
rect 138187 756 138218 8529
rect 138187 752 138252 756
rect 82812 730 138252 752
rect 82812 696 83084 730
rect 138192 696 138252 730
rect 138316 610 138360 8671
rect 82812 523 138360 610
rect 82812 464 83084 523
rect 138307 514 138360 523
rect 138412 8744 138458 8755
rect 138412 524 138424 8744
rect 138458 8182 139132 8216
rect 157792 8182 157852 8216
rect 138458 8156 157852 8182
rect 138458 8019 139072 8156
rect 138458 1278 139072 1414
rect 139106 8094 157818 8156
rect 139106 1340 139189 8094
rect 142463 7594 142510 7660
rect 145055 7594 145102 7660
rect 147638 7594 147702 7660
rect 150228 7594 150292 7660
rect 152822 7594 152886 7660
rect 155412 7594 155476 7660
rect 141509 6766 141679 6782
rect 141509 6664 141525 6766
rect 141658 6664 141679 6766
rect 144101 6766 144271 6782
rect 141509 6648 141679 6664
rect 144101 6664 144117 6766
rect 144250 6664 144271 6766
rect 146693 6766 146863 6782
rect 144101 6648 144271 6664
rect 146693 6664 146709 6766
rect 146842 6664 146863 6766
rect 149269 6766 149455 6782
rect 146693 6648 146863 6664
rect 149269 6664 149301 6766
rect 149434 6664 149455 6766
rect 151877 6766 152047 6782
rect 149269 6648 149455 6664
rect 151877 6664 151893 6766
rect 152026 6664 152047 6766
rect 154469 6766 154639 6782
rect 151877 6648 152047 6664
rect 154469 6664 154485 6766
rect 154618 6664 154639 6766
rect 157061 6766 157231 6782
rect 154469 6648 154639 6664
rect 157061 6664 157077 6766
rect 157210 6664 157231 6766
rect 157061 6648 157231 6664
rect 142463 5966 142510 6032
rect 145055 5966 145102 6032
rect 147638 5966 147702 6032
rect 150228 5966 150292 6032
rect 152818 5966 152882 6032
rect 155416 5966 155480 6032
rect 141509 5138 141679 5154
rect 141509 5036 141525 5138
rect 141658 5036 141679 5138
rect 144101 5138 144271 5154
rect 141509 5020 141679 5036
rect 144101 5036 144117 5138
rect 144250 5036 144271 5138
rect 146677 5138 146863 5154
rect 144101 5020 144271 5036
rect 146677 5036 146709 5138
rect 146842 5036 146863 5138
rect 149285 5138 149455 5154
rect 146677 5020 146863 5036
rect 149285 5036 149301 5138
rect 149434 5036 149455 5138
rect 151877 5138 152047 5154
rect 149285 5020 149455 5036
rect 151877 5036 151893 5138
rect 152026 5036 152047 5138
rect 154469 5138 154639 5154
rect 151877 5020 152047 5036
rect 154469 5036 154485 5138
rect 154618 5036 154639 5138
rect 157061 5138 157231 5154
rect 154469 5020 154639 5036
rect 157061 5036 157077 5138
rect 157210 5036 157231 5138
rect 157061 5020 157231 5036
rect 142463 4338 142510 4404
rect 145055 4338 145102 4404
rect 147638 4338 147702 4404
rect 150226 4338 150290 4404
rect 152822 4338 152886 4404
rect 155414 4338 155478 4404
rect 141509 3510 141679 3526
rect 141509 3408 141525 3510
rect 141658 3408 141679 3510
rect 144101 3510 144271 3526
rect 141509 3392 141679 3408
rect 144101 3408 144117 3510
rect 144250 3408 144271 3510
rect 146693 3510 146863 3526
rect 144101 3392 144271 3408
rect 146693 3408 146709 3510
rect 146842 3408 146863 3510
rect 149285 3510 149455 3526
rect 146693 3392 146863 3408
rect 149285 3408 149301 3510
rect 149434 3408 149455 3510
rect 151877 3510 152047 3526
rect 149285 3392 149455 3408
rect 151877 3408 151893 3510
rect 152026 3408 152047 3510
rect 154469 3510 154639 3526
rect 151877 3392 152047 3408
rect 154469 3408 154485 3510
rect 154618 3408 154639 3510
rect 157061 3510 157231 3526
rect 154469 3392 154639 3408
rect 157061 3408 157077 3510
rect 157210 3408 157231 3510
rect 157061 3392 157231 3408
rect 142463 2710 142510 2776
rect 145055 2710 145102 2776
rect 147638 2710 147702 2776
rect 150226 2710 150290 2776
rect 152642 2770 152926 2776
rect 152642 2716 152664 2770
rect 152900 2716 152926 2770
rect 152642 2710 152926 2716
rect 155416 2710 155480 2776
rect 141509 1882 141679 1898
rect 141509 1780 141525 1882
rect 141658 1780 141679 1882
rect 144101 1882 144271 1898
rect 141509 1764 141679 1780
rect 144101 1780 144117 1882
rect 144250 1780 144271 1882
rect 146693 1882 146863 1898
rect 144101 1764 144271 1780
rect 146693 1780 146709 1882
rect 146842 1780 146863 1882
rect 149285 1882 149455 1898
rect 146693 1764 146863 1780
rect 149285 1780 149301 1882
rect 149434 1780 149455 1882
rect 151877 1882 152047 1898
rect 149285 1764 149455 1780
rect 151877 1780 151893 1882
rect 152026 1780 152047 1882
rect 154469 1882 154639 1898
rect 151877 1764 152047 1780
rect 154469 1780 154485 1882
rect 154618 1780 154639 1882
rect 157061 1882 157231 1898
rect 154469 1764 154639 1780
rect 157061 1780 157077 1882
rect 157210 1780 157231 1882
rect 157061 1764 157231 1780
rect 157724 1340 157818 8094
rect 139106 1278 157818 1340
rect 138458 1252 157852 1278
rect 138458 1218 139132 1252
rect 157792 1218 157852 1252
rect 138458 1217 139161 1218
rect 138412 514 138458 524
rect 138307 498 138458 514
rect 138398 464 138458 498
<< viali >>
rect 137381 8426 137531 8492
rect 138128 752 138187 8529
rect 83084 498 138307 523
rect 138360 514 138412 8755
rect 142129 7624 142175 7803
rect 144721 7624 144767 7803
rect 147313 7624 147359 7803
rect 149905 7624 149951 7803
rect 152497 7624 152543 7803
rect 155089 7624 155135 7803
rect 139918 7316 139966 7547
rect 139782 6677 139816 6781
rect 141525 6664 141658 6766
rect 142374 6677 142408 6781
rect 144117 6664 144250 6766
rect 144966 6677 145000 6781
rect 146709 6664 146842 6766
rect 147558 6677 147592 6781
rect 149301 6664 149434 6766
rect 150150 6677 150184 6781
rect 151893 6664 152026 6766
rect 152742 6677 152776 6781
rect 154485 6664 154618 6766
rect 155334 6677 155368 6781
rect 157077 6664 157210 6766
rect 142129 5996 142175 6175
rect 144721 5996 144767 6175
rect 147313 5996 147359 6175
rect 149905 5996 149951 6175
rect 152497 5996 152543 6175
rect 155089 5996 155135 6175
rect 139918 5688 139966 5919
rect 139782 5049 139816 5153
rect 141525 5036 141658 5138
rect 142374 5049 142408 5153
rect 144117 5036 144250 5138
rect 144966 5049 145000 5153
rect 146709 5036 146842 5138
rect 147558 5049 147592 5153
rect 149301 5036 149434 5138
rect 150150 5049 150184 5153
rect 151893 5036 152026 5138
rect 152742 5049 152776 5153
rect 154485 5036 154618 5138
rect 155334 5049 155368 5153
rect 157077 5036 157210 5138
rect 142129 4368 142175 4547
rect 144721 4368 144767 4547
rect 147313 4368 147359 4547
rect 149905 4368 149951 4547
rect 152497 4368 152543 4547
rect 155089 4368 155135 4547
rect 139918 4060 139966 4291
rect 139782 3421 139816 3525
rect 141525 3408 141658 3510
rect 142374 3421 142408 3525
rect 144117 3408 144250 3510
rect 144966 3421 145000 3525
rect 146709 3408 146842 3510
rect 147558 3421 147592 3525
rect 149301 3408 149434 3510
rect 150150 3421 150184 3525
rect 151893 3408 152026 3510
rect 152742 3421 152776 3525
rect 154485 3408 154618 3510
rect 155334 3421 155368 3525
rect 157077 3408 157210 3510
rect 142129 2740 142175 2919
rect 144721 2740 144767 2919
rect 147313 2740 147359 2919
rect 149905 2740 149951 2919
rect 152497 2740 152543 2919
rect 152664 2716 152900 2770
rect 155089 2740 155135 2919
rect 139918 2432 139966 2663
rect 139782 1793 139816 1897
rect 141525 1780 141658 1882
rect 142374 1793 142408 1897
rect 144117 1780 144250 1882
rect 144966 1793 145000 1897
rect 146709 1780 146842 1882
rect 147558 1793 147592 1897
rect 149301 1780 149434 1882
rect 150150 1793 150184 1897
rect 151893 1780 152026 1882
rect 152742 1793 152776 1897
rect 154485 1780 154618 1882
rect 155334 1793 155368 1897
rect 157077 1780 157210 1882
rect 83084 479 138307 498
<< metal1 >>
rect 138332 8755 138448 8797
rect 103052 8552 103366 8702
rect 103314 7528 103366 8552
rect 106830 8470 106852 8534
rect 138093 8529 138231 8580
rect 137365 8498 137544 8504
rect 138093 8498 138128 8529
rect 137365 8492 138128 8498
rect 137365 8481 137381 8492
rect 137230 8429 137381 8481
rect 137365 8426 137381 8429
rect 137531 8428 138128 8492
rect 137531 8426 137544 8428
rect 137365 8416 137544 8426
rect 138093 6299 138128 8428
rect 138187 6299 138231 8529
rect 138093 4657 138108 6299
rect 138215 4657 138231 6299
rect 84635 1218 84687 1586
rect 137501 1392 137553 1586
rect 137228 1340 137553 1392
rect 84392 1166 84687 1218
rect 138093 752 138128 4657
rect 138187 752 138231 4657
rect 138093 705 138231 752
rect 138332 542 138360 8755
rect 138412 2512 138448 8755
rect 139334 8031 157636 8045
rect 139334 7872 140023 8031
rect 141298 7891 157636 8031
rect 141298 7872 147262 7891
rect 147270 7872 149854 7891
rect 149862 7872 152446 7891
rect 152454 7872 155038 7891
rect 155046 7872 157636 7891
rect 142116 7815 142180 7816
rect 142116 7814 142181 7815
rect 138654 7424 138660 7624
rect 138712 7584 139967 7624
rect 142116 7614 142122 7814
rect 142174 7803 142181 7814
rect 142175 7624 142181 7803
rect 142174 7614 142181 7624
rect 142122 7612 142181 7614
rect 144712 7814 144776 7816
rect 144712 7614 144718 7814
rect 144770 7614 144776 7814
rect 144712 7612 144776 7614
rect 147304 7814 147368 7816
rect 147304 7614 147310 7814
rect 147362 7614 147368 7814
rect 147304 7612 147368 7614
rect 149896 7814 149960 7816
rect 149896 7614 149902 7814
rect 149954 7614 149960 7814
rect 149896 7612 149960 7614
rect 152488 7814 152552 7816
rect 152488 7614 152494 7814
rect 152546 7614 152552 7814
rect 152488 7612 152552 7614
rect 155080 7814 155144 7816
rect 155080 7614 155086 7814
rect 155138 7614 155144 7814
rect 155080 7612 155144 7614
rect 138712 7424 138718 7584
rect 139927 7553 139967 7584
rect 139906 7547 139982 7553
rect 139906 7316 139918 7547
rect 139966 7316 139982 7547
rect 142140 7529 142180 7612
rect 144728 7600 144768 7612
rect 147320 7600 147360 7612
rect 149912 7600 149952 7612
rect 152504 7600 152544 7612
rect 155096 7600 155136 7612
rect 139906 7310 139982 7316
rect 139334 7066 142601 7239
rect 143880 7066 157625 7239
rect 139334 6946 145336 7003
rect 146636 6946 147840 7003
rect 149228 6946 150432 7003
rect 151820 6946 153024 7003
rect 154412 6946 155616 7003
rect 139770 6781 139828 6793
rect 139770 6677 139782 6781
rect 139816 6743 139828 6781
rect 141509 6766 141679 6782
rect 141509 6743 141525 6766
rect 139816 6702 141525 6743
rect 139816 6677 139828 6702
rect 139770 6665 139828 6677
rect 141509 6664 141525 6702
rect 141658 6664 141679 6766
rect 142362 6781 142420 6793
rect 142362 6677 142374 6781
rect 142408 6743 142420 6781
rect 144101 6766 144271 6782
rect 144101 6743 144117 6766
rect 142408 6702 144117 6743
rect 142408 6677 142420 6702
rect 142362 6665 142420 6677
rect 141509 6648 141679 6664
rect 144101 6664 144117 6702
rect 144250 6664 144271 6766
rect 144954 6781 145012 6793
rect 144954 6677 144966 6781
rect 145000 6743 145012 6781
rect 146693 6766 146863 6782
rect 146693 6743 146709 6766
rect 145000 6702 146709 6743
rect 145000 6677 145012 6702
rect 144954 6665 145012 6677
rect 144101 6648 144271 6664
rect 146693 6664 146709 6702
rect 146842 6664 146863 6766
rect 147546 6781 147604 6793
rect 147546 6677 147558 6781
rect 147592 6743 147604 6781
rect 149269 6766 149455 6782
rect 149269 6743 149301 6766
rect 147592 6702 149301 6743
rect 147592 6677 147604 6702
rect 147546 6665 147604 6677
rect 146693 6648 146863 6664
rect 149269 6664 149301 6702
rect 149434 6664 149455 6766
rect 150138 6781 150196 6793
rect 150138 6677 150150 6781
rect 150184 6743 150196 6781
rect 151877 6766 152047 6782
rect 151877 6743 151893 6766
rect 150184 6702 151893 6743
rect 150184 6677 150196 6702
rect 150138 6665 150196 6677
rect 149269 6648 149455 6664
rect 151877 6664 151893 6702
rect 152026 6664 152047 6766
rect 152730 6781 152788 6793
rect 152730 6677 152742 6781
rect 152776 6743 152788 6781
rect 154469 6766 154639 6782
rect 154469 6743 154485 6766
rect 152776 6702 154485 6743
rect 152776 6677 152788 6702
rect 152730 6665 152788 6677
rect 151877 6648 152047 6664
rect 154469 6664 154485 6702
rect 154618 6664 154639 6766
rect 155322 6781 155380 6793
rect 155322 6677 155334 6781
rect 155368 6743 155380 6781
rect 157061 6766 157231 6782
rect 157061 6743 157077 6766
rect 155368 6702 157077 6743
rect 155368 6677 155380 6702
rect 155322 6665 155380 6677
rect 154469 6648 154639 6664
rect 157061 6664 157077 6702
rect 157210 6664 157231 6766
rect 157061 6648 157231 6664
rect 139334 6249 140026 6422
rect 141296 6263 157625 6422
rect 141296 6249 147262 6263
rect 147270 6249 149854 6263
rect 149862 6249 152446 6263
rect 152454 6249 155038 6263
rect 155046 6249 157625 6263
rect 142116 6186 142182 6188
rect 144714 6186 144773 6187
rect 147306 6186 147365 6187
rect 149898 6186 149957 6187
rect 152490 6186 152549 6187
rect 155082 6186 155141 6187
rect 138760 5796 138766 5996
rect 138818 5956 139967 5996
rect 142116 5986 142122 6186
rect 142174 6175 142182 6186
rect 142175 5996 142182 6175
rect 142174 5986 142182 5996
rect 144712 5986 144718 6186
rect 144770 5986 144776 6186
rect 142122 5984 142181 5986
rect 144712 5984 144776 5986
rect 147304 5986 147310 6186
rect 147362 5986 147368 6186
rect 147304 5984 147368 5986
rect 149896 5986 149902 6186
rect 149954 5986 149960 6186
rect 149896 5984 149960 5986
rect 152488 5986 152494 6186
rect 152546 5986 152552 6186
rect 152488 5984 152552 5986
rect 155080 5986 155086 6186
rect 155138 5986 155144 6186
rect 155080 5984 155144 5986
rect 138818 5796 138824 5956
rect 139927 5925 139967 5956
rect 139906 5919 139982 5925
rect 139906 5688 139918 5919
rect 139966 5688 139982 5919
rect 142140 5901 142180 5984
rect 144728 5980 144768 5984
rect 147320 5980 147360 5984
rect 149912 5980 149952 5984
rect 152504 5980 152544 5984
rect 155096 5980 155136 5984
rect 139906 5682 139982 5688
rect 139334 5438 142597 5611
rect 143876 5438 157642 5611
rect 139334 5318 145336 5375
rect 146636 5318 147840 5375
rect 149228 5318 150432 5375
rect 151820 5318 153024 5375
rect 154412 5318 155616 5375
rect 139770 5153 139828 5165
rect 139770 5049 139782 5153
rect 139816 5115 139828 5153
rect 141509 5138 141679 5154
rect 141509 5115 141525 5138
rect 139816 5074 141525 5115
rect 139816 5049 139828 5074
rect 139770 5037 139828 5049
rect 141509 5036 141525 5074
rect 141658 5036 141679 5138
rect 142362 5153 142420 5165
rect 142362 5049 142374 5153
rect 142408 5115 142420 5153
rect 144101 5138 144271 5154
rect 144101 5115 144117 5138
rect 142408 5074 144117 5115
rect 142408 5049 142420 5074
rect 142362 5037 142420 5049
rect 141509 5020 141679 5036
rect 144101 5036 144117 5074
rect 144250 5036 144271 5138
rect 144954 5153 145012 5165
rect 144954 5049 144966 5153
rect 145000 5115 145012 5153
rect 146677 5138 146863 5154
rect 146677 5115 146709 5138
rect 145000 5074 146709 5115
rect 145000 5049 145012 5074
rect 144954 5037 145012 5049
rect 144101 5020 144271 5036
rect 146677 5036 146709 5074
rect 146842 5036 146863 5138
rect 147546 5153 147604 5165
rect 147546 5049 147558 5153
rect 147592 5115 147604 5153
rect 149285 5138 149455 5154
rect 149285 5115 149301 5138
rect 147592 5074 149301 5115
rect 147592 5049 147604 5074
rect 147546 5037 147604 5049
rect 146677 5020 146863 5036
rect 149285 5036 149301 5074
rect 149434 5036 149455 5138
rect 150138 5153 150196 5165
rect 150138 5049 150150 5153
rect 150184 5115 150196 5153
rect 151877 5138 152047 5154
rect 151877 5115 151893 5138
rect 150184 5074 151893 5115
rect 150184 5049 150196 5074
rect 150138 5037 150196 5049
rect 149285 5020 149455 5036
rect 151877 5036 151893 5074
rect 152026 5036 152047 5138
rect 152730 5153 152788 5165
rect 152730 5049 152742 5153
rect 152776 5115 152788 5153
rect 154469 5138 154639 5154
rect 154469 5115 154485 5138
rect 152776 5074 154485 5115
rect 152776 5049 152788 5074
rect 152730 5037 152788 5049
rect 151877 5020 152047 5036
rect 154469 5036 154485 5074
rect 154618 5036 154639 5138
rect 155322 5153 155380 5165
rect 155322 5049 155334 5153
rect 155368 5115 155380 5153
rect 157061 5138 157231 5154
rect 157061 5115 157077 5138
rect 155368 5074 157077 5115
rect 155368 5049 155380 5074
rect 155322 5037 155380 5049
rect 154469 5020 154639 5036
rect 157061 5036 157077 5074
rect 157210 5036 157231 5138
rect 157061 5020 157231 5036
rect 139334 4622 140024 4795
rect 141294 4731 157614 4795
rect 141294 4697 147319 4731
rect 147353 4697 149911 4731
rect 149945 4706 152503 4731
rect 149945 4697 150007 4706
rect 150014 4697 152503 4706
rect 152537 4706 155095 4731
rect 152537 4697 152599 4706
rect 152606 4697 155095 4706
rect 155129 4706 157614 4731
rect 155129 4697 155191 4706
rect 155198 4697 157614 4706
rect 141294 4635 157614 4697
rect 141294 4622 147266 4635
rect 147270 4622 149858 4635
rect 149862 4622 152450 4635
rect 152454 4622 155042 4635
rect 155046 4622 157614 4635
rect 142116 4559 142180 4560
rect 142116 4558 142181 4559
rect 144714 4558 144773 4559
rect 147306 4558 147365 4559
rect 149898 4558 149957 4559
rect 152490 4558 152549 4559
rect 155082 4558 155141 4559
rect 142116 4528 142122 4558
rect 142174 4547 142181 4558
rect 138842 4168 138848 4368
rect 138900 4328 139967 4368
rect 142116 4358 142122 4488
rect 142175 4368 142181 4547
rect 142174 4358 142181 4368
rect 142122 4356 142181 4358
rect 144712 4358 144718 4558
rect 144770 4358 144776 4558
rect 144712 4356 144776 4358
rect 147304 4358 147310 4558
rect 147362 4358 147368 4558
rect 147304 4356 147368 4358
rect 149896 4358 149902 4558
rect 149954 4358 149960 4558
rect 149896 4356 149960 4358
rect 152488 4358 152494 4558
rect 152546 4358 152552 4558
rect 152488 4356 152552 4358
rect 155080 4358 155086 4558
rect 155138 4358 155144 4558
rect 155080 4356 155144 4358
rect 144728 4350 144768 4356
rect 147320 4350 147360 4356
rect 149912 4350 149952 4356
rect 152504 4350 152544 4356
rect 155096 4350 155136 4356
rect 138900 4168 138906 4328
rect 139927 4297 139967 4328
rect 139906 4291 139982 4297
rect 139906 4060 139918 4291
rect 139966 4060 139982 4291
rect 139906 4054 139982 4060
rect 139334 3822 142601 3995
rect 143880 3822 157631 3995
rect 139334 3690 145336 3747
rect 146636 3690 147840 3747
rect 149228 3690 150432 3747
rect 151820 3690 153024 3747
rect 154412 3690 155616 3747
rect 139770 3525 139828 3537
rect 139770 3421 139782 3525
rect 139816 3487 139828 3525
rect 141509 3510 141679 3526
rect 141509 3487 141525 3510
rect 139816 3446 141525 3487
rect 139816 3421 139828 3446
rect 139770 3409 139828 3421
rect 141509 3408 141525 3446
rect 141658 3408 141679 3510
rect 142362 3525 142420 3537
rect 142362 3421 142374 3525
rect 142408 3487 142420 3525
rect 144101 3510 144271 3526
rect 144101 3487 144117 3510
rect 142408 3446 144117 3487
rect 142408 3421 142420 3446
rect 142362 3409 142420 3421
rect 141509 3392 141679 3408
rect 144101 3408 144117 3446
rect 144250 3408 144271 3510
rect 144954 3525 145012 3537
rect 144954 3421 144966 3525
rect 145000 3487 145012 3525
rect 146693 3510 146863 3526
rect 146693 3487 146709 3510
rect 145000 3446 146709 3487
rect 145000 3421 145012 3446
rect 144954 3409 145012 3421
rect 144101 3392 144271 3408
rect 146693 3408 146709 3446
rect 146842 3408 146863 3510
rect 147546 3525 147604 3537
rect 147546 3421 147558 3525
rect 147592 3487 147604 3525
rect 149285 3510 149455 3526
rect 149285 3487 149301 3510
rect 147592 3446 149301 3487
rect 147592 3421 147604 3446
rect 147546 3409 147604 3421
rect 146693 3392 146863 3408
rect 149285 3408 149301 3446
rect 149434 3408 149455 3510
rect 150138 3525 150196 3537
rect 150138 3421 150150 3525
rect 150184 3487 150196 3525
rect 151877 3510 152047 3526
rect 151877 3487 151893 3510
rect 150184 3446 151893 3487
rect 150184 3421 150196 3446
rect 150138 3409 150196 3421
rect 149285 3392 149455 3408
rect 151877 3408 151893 3446
rect 152026 3408 152047 3510
rect 152730 3525 152788 3537
rect 152730 3421 152742 3525
rect 152776 3487 152788 3525
rect 154469 3510 154639 3526
rect 154469 3487 154485 3510
rect 152776 3446 154485 3487
rect 152776 3421 152788 3446
rect 152730 3409 152788 3421
rect 151877 3392 152047 3408
rect 154469 3408 154485 3446
rect 154618 3408 154639 3510
rect 155322 3525 155380 3537
rect 155322 3421 155334 3525
rect 155368 3487 155380 3525
rect 157061 3510 157231 3526
rect 157061 3487 157077 3510
rect 155368 3446 157077 3487
rect 155368 3421 155380 3446
rect 155322 3409 155380 3421
rect 154469 3392 154639 3408
rect 157061 3408 157077 3446
rect 157210 3408 157231 3510
rect 157061 3392 157231 3408
rect 138932 2828 138938 3028
rect 138990 2869 138996 3028
rect 139334 3000 140028 3173
rect 141298 3007 157598 3173
rect 141298 3000 147252 3007
rect 147270 3000 149844 3007
rect 149862 3000 152436 3007
rect 152454 3000 155028 3007
rect 155046 3000 157598 3007
rect 142116 2930 142182 2932
rect 144714 2930 144773 2931
rect 147306 2930 147365 2931
rect 149898 2930 149957 2931
rect 152490 2930 152549 2931
rect 155082 2930 155141 2931
rect 142116 2900 142122 2930
rect 142174 2919 142182 2930
rect 138990 2828 140215 2869
rect 138981 2827 140215 2828
rect 139032 2540 139038 2740
rect 139090 2700 139963 2740
rect 139090 2540 139096 2700
rect 139923 2669 139963 2700
rect 139906 2663 139979 2669
rect 138412 2481 138622 2512
rect 138593 1342 138622 2481
rect 139906 2432 139918 2663
rect 139966 2432 139979 2663
rect 140173 2558 140215 2827
rect 142116 2730 142122 2860
rect 142175 2740 142182 2919
rect 142174 2730 142182 2740
rect 144712 2730 144718 2930
rect 144770 2730 144776 2930
rect 142122 2728 142181 2730
rect 144712 2728 144776 2730
rect 147304 2730 147310 2930
rect 147362 2730 147368 2930
rect 147304 2728 147368 2730
rect 149896 2730 149902 2930
rect 149954 2730 149960 2930
rect 149896 2728 149960 2730
rect 152488 2730 152494 2930
rect 152546 2730 152552 2930
rect 152488 2728 152552 2730
rect 152642 2770 152926 2776
rect 144728 2710 144768 2728
rect 147320 2710 147360 2728
rect 149912 2710 149952 2728
rect 152504 2710 152544 2728
rect 152642 2716 152664 2770
rect 152900 2716 152926 2770
rect 155080 2730 155086 2930
rect 155138 2730 155144 2930
rect 155080 2728 155144 2730
rect 152642 2710 152926 2716
rect 155096 2710 155136 2728
rect 152681 2558 152723 2710
rect 140173 2516 152723 2558
rect 139906 2426 139979 2432
rect 139334 2183 142601 2356
rect 143880 2183 157642 2356
rect 139334 2062 145336 2119
rect 146636 2062 147840 2119
rect 149228 2062 150432 2119
rect 151820 2062 153024 2119
rect 154412 2062 155616 2119
rect 139770 1897 139828 1909
rect 139770 1793 139782 1897
rect 139816 1859 139828 1897
rect 141509 1882 141679 1898
rect 141509 1859 141525 1882
rect 139816 1818 141525 1859
rect 139816 1793 139828 1818
rect 139770 1781 139828 1793
rect 141509 1780 141525 1818
rect 141658 1780 141679 1882
rect 142362 1897 142420 1909
rect 142362 1793 142374 1897
rect 142408 1859 142420 1897
rect 144101 1882 144271 1898
rect 144101 1859 144117 1882
rect 142408 1818 144117 1859
rect 142408 1793 142420 1818
rect 142362 1781 142420 1793
rect 141509 1764 141679 1780
rect 144101 1780 144117 1818
rect 144250 1780 144271 1882
rect 144954 1897 145012 1909
rect 144954 1793 144966 1897
rect 145000 1859 145012 1897
rect 146693 1882 146863 1898
rect 146693 1859 146709 1882
rect 145000 1818 146709 1859
rect 145000 1793 145012 1818
rect 144954 1781 145012 1793
rect 144101 1764 144271 1780
rect 146693 1780 146709 1818
rect 146842 1780 146863 1882
rect 147546 1897 147604 1909
rect 147546 1793 147558 1897
rect 147592 1859 147604 1897
rect 149285 1882 149455 1898
rect 149285 1859 149301 1882
rect 147592 1818 149301 1859
rect 147592 1793 147604 1818
rect 147546 1781 147604 1793
rect 146693 1764 146863 1780
rect 149285 1780 149301 1818
rect 149434 1780 149455 1882
rect 150138 1897 150196 1909
rect 150138 1793 150150 1897
rect 150184 1859 150196 1897
rect 151877 1882 152047 1898
rect 151877 1859 151893 1882
rect 150184 1818 151893 1859
rect 150184 1793 150196 1818
rect 150138 1781 150196 1793
rect 149285 1764 149455 1780
rect 151877 1780 151893 1818
rect 152026 1780 152047 1882
rect 152730 1897 152788 1909
rect 152730 1793 152742 1897
rect 152776 1859 152788 1897
rect 154469 1882 154639 1898
rect 154469 1859 154485 1882
rect 152776 1818 154485 1859
rect 152776 1793 152788 1818
rect 152730 1781 152788 1793
rect 151877 1764 152047 1780
rect 154469 1780 154485 1818
rect 154618 1780 154639 1882
rect 155322 1897 155380 1909
rect 155322 1793 155334 1897
rect 155368 1859 155380 1897
rect 157061 1882 157231 1898
rect 157061 1859 157077 1882
rect 155368 1818 157077 1859
rect 155368 1793 155380 1818
rect 155322 1781 155380 1793
rect 154469 1764 154639 1780
rect 157061 1780 157077 1818
rect 157210 1780 157231 1882
rect 157061 1764 157231 1780
rect 139334 1461 140021 1539
rect 141293 1461 157564 1539
rect 82812 523 138360 542
rect 82812 479 83084 523
rect 138307 514 138360 523
rect 138412 1310 138622 1342
rect 138412 514 138448 1310
rect 138307 479 138448 514
rect 82812 464 138448 479
<< via1 >>
rect 138108 4657 138128 6299
rect 138128 4657 138187 6299
rect 138187 4657 138215 6299
rect 140023 7868 141298 8031
rect 138660 7424 138712 7624
rect 142122 7803 142174 7814
rect 142122 7624 142129 7803
rect 142129 7624 142174 7803
rect 142122 7614 142174 7624
rect 144718 7803 144770 7814
rect 144718 7624 144721 7803
rect 144721 7624 144767 7803
rect 144767 7624 144770 7803
rect 144718 7614 144770 7624
rect 147310 7803 147362 7814
rect 147310 7624 147313 7803
rect 147313 7624 147359 7803
rect 147359 7624 147362 7803
rect 147310 7614 147362 7624
rect 149902 7803 149954 7814
rect 149902 7624 149905 7803
rect 149905 7624 149951 7803
rect 149951 7624 149954 7803
rect 149902 7614 149954 7624
rect 152494 7803 152546 7814
rect 152494 7624 152497 7803
rect 152497 7624 152543 7803
rect 152543 7624 152546 7803
rect 152494 7614 152546 7624
rect 155086 7803 155138 7814
rect 155086 7624 155089 7803
rect 155089 7624 155135 7803
rect 155135 7624 155138 7803
rect 155086 7614 155138 7624
rect 142601 7047 143880 7264
rect 145336 6946 146330 7003
rect 141525 6664 141658 6766
rect 144117 6664 144250 6766
rect 146709 6664 146842 6766
rect 149301 6664 149434 6766
rect 151893 6664 152026 6766
rect 154485 6664 154618 6766
rect 157077 6664 157210 6766
rect 140026 6229 141296 6444
rect 138766 5796 138818 5996
rect 142122 6175 142174 6186
rect 142122 5996 142129 6175
rect 142129 5996 142174 6175
rect 142122 5986 142174 5996
rect 144718 6175 144770 6186
rect 144718 5996 144721 6175
rect 144721 5996 144767 6175
rect 144767 5996 144770 6175
rect 144718 5986 144770 5996
rect 147310 6175 147362 6186
rect 147310 5996 147313 6175
rect 147313 5996 147359 6175
rect 147359 5996 147362 6175
rect 147310 5986 147362 5996
rect 149902 6175 149954 6186
rect 149902 5996 149905 6175
rect 149905 5996 149951 6175
rect 149951 5996 149954 6175
rect 149902 5986 149954 5996
rect 152494 6175 152546 6186
rect 152494 5996 152497 6175
rect 152497 5996 152543 6175
rect 152543 5996 152546 6175
rect 152494 5986 152546 5996
rect 155086 6175 155138 6186
rect 155086 5996 155089 6175
rect 155089 5996 155135 6175
rect 155135 5996 155138 6175
rect 155086 5986 155138 5996
rect 142597 5420 143876 5637
rect 145336 5318 146330 5375
rect 141525 5036 141658 5138
rect 144117 5036 144250 5138
rect 146709 5036 146842 5138
rect 149301 5036 149434 5138
rect 151893 5036 152026 5138
rect 154485 5036 154618 5138
rect 157077 5036 157210 5138
rect 140024 4609 141294 4824
rect 142122 4547 142174 4558
rect 138848 4168 138900 4368
rect 142122 4368 142129 4547
rect 142129 4368 142174 4547
rect 142122 4358 142174 4368
rect 144718 4547 144770 4558
rect 144718 4368 144721 4547
rect 144721 4368 144767 4547
rect 144767 4368 144770 4547
rect 144718 4358 144770 4368
rect 147310 4547 147362 4558
rect 147310 4368 147313 4547
rect 147313 4368 147359 4547
rect 147359 4368 147362 4547
rect 147310 4358 147362 4368
rect 149902 4547 149954 4558
rect 149902 4368 149905 4547
rect 149905 4368 149951 4547
rect 149951 4368 149954 4547
rect 149902 4358 149954 4368
rect 152494 4547 152546 4558
rect 152494 4368 152497 4547
rect 152497 4368 152543 4547
rect 152543 4368 152546 4547
rect 152494 4358 152546 4368
rect 155086 4547 155138 4558
rect 155086 4368 155089 4547
rect 155089 4368 155135 4547
rect 155135 4368 155138 4547
rect 155086 4358 155138 4368
rect 142601 3789 143880 4006
rect 145336 3690 146330 3747
rect 141525 3408 141658 3510
rect 144117 3408 144250 3510
rect 146709 3408 146842 3510
rect 149301 3408 149434 3510
rect 151893 3408 152026 3510
rect 154485 3408 154618 3510
rect 157077 3408 157210 3510
rect 138938 2828 138990 3028
rect 140028 2976 141298 3191
rect 142122 2919 142174 2930
rect 139038 2540 139090 2740
rect 138379 1342 138412 2481
rect 138412 1342 138593 2481
rect 142122 2740 142129 2919
rect 142129 2740 142174 2919
rect 142122 2730 142174 2740
rect 144718 2919 144770 2930
rect 144718 2740 144721 2919
rect 144721 2740 144767 2919
rect 144767 2740 144770 2919
rect 144718 2730 144770 2740
rect 147310 2919 147362 2930
rect 147310 2740 147313 2919
rect 147313 2740 147359 2919
rect 147359 2740 147362 2919
rect 147310 2730 147362 2740
rect 149902 2919 149954 2930
rect 149902 2740 149905 2919
rect 149905 2740 149951 2919
rect 149951 2740 149954 2919
rect 149902 2730 149954 2740
rect 152494 2919 152546 2930
rect 152494 2740 152497 2919
rect 152497 2740 152543 2919
rect 152543 2740 152546 2919
rect 152494 2730 152546 2740
rect 155086 2919 155138 2930
rect 155086 2740 155089 2919
rect 155089 2740 155135 2919
rect 155135 2740 155138 2919
rect 155086 2730 155138 2740
rect 142601 2163 143880 2380
rect 145336 2062 146330 2119
rect 141525 1780 141658 1882
rect 144117 1780 144250 1882
rect 146709 1780 146842 1882
rect 149301 1780 149434 1882
rect 151893 1780 152026 1882
rect 154485 1780 154618 1882
rect 157077 1780 157210 1882
rect 140021 1448 141293 1563
<< metal2 >>
rect 93490 11266 155452 11314
rect 83080 8465 92448 8697
rect 92775 8465 93336 8697
rect 93490 8390 93538 11266
rect 103234 11170 155266 11218
rect 93778 8465 102964 8697
rect 83240 8158 93538 8390
rect 93924 8158 103136 8390
rect 103234 8310 103282 11170
rect 104706 11074 155132 11122
rect 103354 8465 103368 8697
rect 103695 8465 104546 8697
rect 104706 8390 104754 11074
rect 106804 10978 154996 11026
rect 104988 8465 105264 8697
rect 105591 8465 106702 8697
rect 106804 8390 106852 10978
rect 112201 10882 152860 10930
rect 107126 8465 111138 8697
rect 111465 8465 112026 8697
rect 112201 8390 112249 10882
rect 103568 8310 103672 8390
rect 103234 8262 103672 8310
rect 103568 8158 103672 8262
rect 104090 8162 104754 8390
rect 104090 8158 104724 8162
rect 105168 8158 106859 8390
rect 107293 8162 112249 8390
rect 112358 10786 152674 10834
rect 112358 8366 112406 10786
rect 114215 10690 152540 10738
rect 112456 8465 113274 8697
rect 113601 8465 114172 8697
rect 114215 8390 114263 10690
rect 114857 10594 152404 10642
rect 114332 8465 114342 8697
rect 114669 8465 114693 8697
rect 114857 8390 114905 10594
rect 121263 10498 150268 10546
rect 115132 8465 120750 8697
rect 121077 8465 121102 8697
rect 121263 8390 121311 10498
rect 112559 8366 112737 8390
rect 112358 8318 112737 8366
rect 107293 8158 112208 8162
rect 112559 8158 112737 8318
rect 113174 8158 114343 8390
rect 114781 8160 114905 8390
rect 115319 8162 121311 8390
rect 121452 10402 150082 10450
rect 121452 8366 121500 10402
rect 126066 10306 149948 10354
rect 121543 8465 125556 8697
rect 125883 8465 125914 8697
rect 126066 8390 126114 10306
rect 121630 8366 121831 8390
rect 121452 8318 121831 8366
rect 114781 8158 114880 8160
rect 115319 8158 121275 8162
rect 121630 8158 121831 8318
rect 122256 8162 126114 8390
rect 126243 10210 149812 10258
rect 126243 8390 126291 10210
rect 127688 10114 147676 10162
rect 126351 8465 127158 8697
rect 127485 8465 127508 8697
rect 127688 8390 127736 10114
rect 126243 8342 126627 8390
rect 122256 8158 126094 8162
rect 126442 8158 126627 8342
rect 127066 8161 127736 8390
rect 127864 10018 147490 10066
rect 127864 8371 127912 10018
rect 129296 9922 147356 9970
rect 127945 8465 128760 8697
rect 129087 8465 129125 8697
rect 129296 8390 129344 9922
rect 128040 8371 128250 8390
rect 127864 8323 128250 8371
rect 127066 8158 127694 8161
rect 128040 8158 128250 8323
rect 128655 8159 129344 8390
rect 129433 9826 147220 9874
rect 129433 8361 129481 9826
rect 130876 9730 145084 9778
rect 129546 8465 130362 8697
rect 130689 8465 130721 8697
rect 130876 8390 130924 9730
rect 129617 8361 129830 8390
rect 129433 8313 129830 8361
rect 128655 8158 129305 8159
rect 129617 8158 129830 8313
rect 130266 8160 130924 8390
rect 131034 9634 144898 9682
rect 131034 8370 131082 9634
rect 132491 9538 144764 9586
rect 131147 8465 131964 8697
rect 132291 8465 132328 8697
rect 132491 8390 132539 9538
rect 131242 8370 131420 8390
rect 131034 8322 131420 8370
rect 130266 8158 130900 8160
rect 131242 8158 131420 8322
rect 131865 8161 132539 8390
rect 132679 9442 144628 9490
rect 132679 8379 132727 9442
rect 134079 9346 142486 9394
rect 132825 8465 133566 8697
rect 133893 8465 133926 8697
rect 134079 8390 134127 9346
rect 132825 8379 133034 8390
rect 132679 8331 133034 8379
rect 131865 8158 132499 8161
rect 132825 8158 133034 8331
rect 133461 8158 134127 8390
rect 134215 9250 142330 9298
rect 134215 8374 134263 9250
rect 135729 9154 142168 9202
rect 134356 8464 134908 8697
rect 134929 8465 135168 8697
rect 135495 8465 135568 8697
rect 135729 8390 135777 9154
rect 134544 8374 134639 8390
rect 134215 8326 134639 8374
rect 134544 8158 134639 8326
rect 135033 8333 135777 8390
rect 135885 9058 142020 9106
rect 135885 8373 135933 9058
rect 135981 8465 135997 8697
rect 136169 8465 136203 8697
rect 136506 8465 137113 8697
rect 135981 8373 136549 8390
rect 135033 8158 135718 8333
rect 135885 8325 136549 8373
rect 135981 8158 136549 8325
rect 136693 8158 137292 8390
rect 140008 8031 141311 8086
rect 82836 7757 137616 7995
rect 140008 7868 140023 8031
rect 141298 7868 141311 8031
rect 82836 7756 82958 7757
rect 137608 7426 137655 7660
rect 137910 7426 137939 7660
rect 138660 7624 138712 7632
rect 138660 7418 138712 7424
rect 82836 6533 137616 6766
rect 83018 6532 137616 6533
rect 138079 6299 138270 6322
rect 82892 5635 137616 5869
rect 82883 4654 83084 4738
rect 137608 4712 137654 4872
rect 137146 4654 137654 4712
rect 137608 4638 137654 4654
rect 137909 4638 137938 4872
rect 138079 4657 138108 6299
rect 138215 4657 138270 6299
rect 138079 4638 138270 4657
rect 82836 4463 108079 4480
rect 82836 4379 83084 4463
rect 82836 4377 83162 4379
rect 82836 4242 108079 4377
rect 82892 3263 137597 3501
rect 138358 2481 138622 2512
rect 82836 1496 137597 1734
rect 138358 1342 138379 2481
rect 138593 1342 138622 2481
rect 138358 1310 138622 1342
rect 135140 1287 135180 1289
rect 83275 1099 90318 1287
rect 90748 1099 130376 1287
rect 130778 1286 133033 1287
rect 130778 1099 133047 1286
rect 133472 1099 134103 1287
rect 134542 1099 135180 1287
rect 135611 1284 136210 1287
rect 135611 1099 136229 1284
rect 136690 1099 137068 1287
rect 137185 1099 137300 1287
rect 83112 843 90152 1031
rect 90582 843 129222 1031
rect 129549 843 130220 1031
rect 130336 152 130376 1099
rect 130622 843 132450 1031
rect 132777 843 132870 1031
rect 133007 240 133047 1099
rect 133309 843 133529 1031
rect 133856 843 133946 1031
rect 134062 330 134102 1099
rect 134385 843 134534 1031
rect 134861 843 135007 1031
rect 135140 412 135180 1099
rect 135446 843 135582 1031
rect 135909 843 136081 1031
rect 136189 518 136229 1099
rect 136525 843 137135 1031
rect 138666 518 138706 7418
rect 139402 7344 139532 7384
rect 140008 6444 141311 7868
rect 141980 7194 142020 9058
rect 142128 7824 142168 9154
rect 142122 7814 142174 7824
rect 142122 7606 142174 7614
rect 141980 7154 142168 7194
rect 141509 6766 141679 6782
rect 141509 6664 141525 6766
rect 141658 6739 141679 6766
rect 141658 6699 142039 6739
rect 141658 6664 141679 6699
rect 141509 6648 141679 6664
rect 140008 6229 140026 6444
rect 141296 6229 141311 6444
rect 138766 5996 138818 6004
rect 138766 5790 138818 5796
rect 136189 478 138706 518
rect 138772 412 138812 5790
rect 140008 4824 141311 6229
rect 141509 5138 141679 5154
rect 141509 5036 141525 5138
rect 141658 5097 141679 5138
rect 141658 5057 141919 5097
rect 141658 5036 141679 5057
rect 141509 5020 141679 5036
rect 140008 4609 140024 4824
rect 141294 4609 141311 4824
rect 138848 4368 138900 4376
rect 138848 4162 138900 4168
rect 135140 372 138812 412
rect 138854 330 138894 4162
rect 140008 3191 141311 4609
rect 141509 3510 141679 3526
rect 141509 3408 141525 3510
rect 141658 3474 141679 3510
rect 141658 3434 141803 3474
rect 141658 3408 141679 3434
rect 141509 3392 141679 3408
rect 138944 3034 138984 3044
rect 138938 3028 138990 3034
rect 138938 2820 138990 2828
rect 140008 2976 140028 3191
rect 141298 2976 141311 3191
rect 134062 290 138894 330
rect 138942 240 138982 2820
rect 139038 2740 139090 2748
rect 139038 2534 139090 2540
rect 133007 200 138982 240
rect 139044 152 139084 2534
rect 140008 2485 141311 2976
rect 140008 1563 140035 2485
rect 141277 1563 141311 2485
rect 141509 1882 141679 1898
rect 141509 1780 141525 1882
rect 141658 1780 141679 1882
rect 141509 1764 141679 1780
rect 140008 1448 140021 1563
rect 141293 1448 141311 1563
rect 140008 1340 140035 1448
rect 141277 1340 141311 1448
rect 140008 1300 141311 1340
rect 141639 678 141679 1764
rect 141759 1096 141803 3434
rect 141763 678 141803 1096
rect 141879 678 141919 5057
rect 141999 678 142039 6699
rect 142128 6196 142168 7154
rect 142122 6186 142174 6196
rect 142122 5978 142174 5986
rect 142290 5302 142330 9250
rect 142128 5262 142330 5302
rect 142128 4568 142168 5262
rect 142122 4558 142174 4568
rect 142122 4350 142174 4358
rect 142446 4076 142486 9346
rect 142128 4036 142486 4076
rect 142588 7264 143893 8101
rect 142588 7047 142601 7264
rect 143880 7047 143893 7264
rect 144588 7178 144628 9442
rect 144724 7824 144764 9538
rect 144718 7814 144770 7824
rect 144718 7606 144770 7614
rect 144588 7138 144764 7178
rect 142588 6280 143893 7047
rect 144101 6766 144271 6782
rect 144101 6664 144117 6766
rect 144250 6739 144271 6766
rect 144250 6699 144631 6739
rect 144250 6664 144271 6699
rect 144101 6648 144271 6664
rect 142588 5637 142647 6280
rect 143849 5637 143893 6280
rect 142588 5420 142597 5637
rect 143876 5420 143893 5637
rect 142588 4689 142647 5420
rect 143849 4689 143893 5420
rect 144101 5138 144271 5154
rect 144101 5036 144117 5138
rect 144250 5097 144271 5138
rect 144250 5057 144511 5097
rect 144250 5036 144271 5057
rect 144101 5020 144271 5036
rect 142128 2940 142168 4036
rect 142588 4006 143893 4689
rect 142588 3789 142601 4006
rect 143880 3789 143893 4006
rect 142122 2930 142174 2940
rect 142122 2722 142174 2730
rect 142588 2380 143893 3789
rect 144101 3510 144271 3526
rect 144101 3408 144117 3510
rect 144250 3474 144271 3510
rect 144250 3434 144391 3474
rect 144250 3408 144271 3434
rect 144101 3392 144271 3408
rect 142588 2163 142601 2380
rect 143880 2163 143893 2380
rect 142588 1390 143893 2163
rect 144101 1882 144271 1898
rect 144101 1780 144117 1882
rect 144250 1780 144271 1882
rect 144101 1764 144271 1780
rect 144231 678 144271 1764
rect 144351 678 144391 3434
rect 144471 678 144511 5057
rect 144591 678 144631 6699
rect 144724 6196 144764 7138
rect 144718 6186 144770 6196
rect 144718 5978 144770 5986
rect 144858 5870 144898 9634
rect 144724 5830 144898 5870
rect 144724 4568 144764 5830
rect 144718 4558 144770 4568
rect 144718 4350 144770 4358
rect 145044 4090 145084 9730
rect 144724 4050 145084 4090
rect 145336 7851 146330 8094
rect 145336 7003 145367 7851
rect 146299 7003 146330 7851
rect 147180 7178 147220 9826
rect 147316 7824 147356 9922
rect 147310 7814 147362 7824
rect 147310 7606 147362 7614
rect 147180 7138 147356 7178
rect 145336 6713 145367 6946
rect 146299 6713 146330 6946
rect 145336 5375 146330 6713
rect 146693 6766 146863 6782
rect 146693 6664 146709 6766
rect 146842 6739 146863 6766
rect 146842 6699 147223 6739
rect 146842 6664 146863 6699
rect 146693 6648 146863 6664
rect 144724 2940 144764 4050
rect 145336 3747 146330 5318
rect 146693 5138 146863 5154
rect 146693 5036 146709 5138
rect 146842 5097 146863 5138
rect 146842 5057 147103 5097
rect 146842 5036 146863 5057
rect 146693 5020 146863 5036
rect 144718 2930 144770 2940
rect 144718 2722 144770 2730
rect 145336 2119 146330 3690
rect 146693 3510 146863 3526
rect 146693 3408 146709 3510
rect 146842 3474 146863 3510
rect 146842 3434 146983 3474
rect 146842 3408 146863 3434
rect 146693 3392 146863 3408
rect 145336 1301 146330 2062
rect 146693 1882 146863 1898
rect 146693 1780 146709 1882
rect 146842 1780 146863 1882
rect 146693 1764 146863 1780
rect 146823 678 146863 1764
rect 146943 678 146983 3434
rect 147063 678 147103 5057
rect 147183 678 147223 6699
rect 147316 6196 147356 7138
rect 147310 6186 147362 6196
rect 147310 5978 147362 5986
rect 147450 5870 147490 10018
rect 147316 5830 147490 5870
rect 147316 4568 147356 5830
rect 147310 4558 147362 4568
rect 147310 4350 147362 4358
rect 147636 4090 147676 10114
rect 149772 7178 149812 10210
rect 149908 7824 149948 10306
rect 149902 7814 149954 7824
rect 149902 7606 149954 7614
rect 149772 7138 149948 7178
rect 149285 6766 149455 6782
rect 149285 6664 149301 6766
rect 149434 6739 149455 6766
rect 149434 6699 149815 6739
rect 149434 6664 149455 6699
rect 149285 6648 149455 6664
rect 149285 5138 149455 5154
rect 149285 5036 149301 5138
rect 149434 5097 149455 5138
rect 149434 5057 149695 5097
rect 149434 5036 149455 5057
rect 149285 5020 149455 5036
rect 147316 4050 147676 4090
rect 147316 2940 147356 4050
rect 149285 3510 149455 3526
rect 149285 3408 149301 3510
rect 149434 3474 149455 3510
rect 149434 3434 149575 3474
rect 149434 3408 149455 3434
rect 149285 3392 149455 3408
rect 147310 2930 147362 2940
rect 147310 2722 147362 2730
rect 149285 1882 149455 1898
rect 149285 1780 149301 1882
rect 149434 1780 149455 1882
rect 149285 1764 149455 1780
rect 149415 678 149455 1764
rect 149535 678 149575 3434
rect 149655 678 149695 5057
rect 149775 678 149815 6699
rect 149908 6196 149948 7138
rect 149902 6186 149954 6196
rect 149902 5978 149954 5986
rect 150042 5870 150082 10402
rect 149908 5830 150082 5870
rect 149908 4568 149948 5830
rect 149902 4558 149954 4568
rect 149902 4350 149954 4358
rect 150228 4090 150268 10498
rect 152364 7178 152404 10594
rect 152500 7824 152540 10690
rect 152494 7814 152546 7824
rect 152494 7606 152546 7614
rect 152364 7138 152540 7178
rect 151877 6766 152047 6782
rect 151877 6664 151893 6766
rect 152026 6739 152047 6766
rect 152026 6699 152407 6739
rect 152026 6664 152047 6699
rect 151877 6648 152047 6664
rect 151877 5138 152047 5154
rect 151877 5036 151893 5138
rect 152026 5097 152047 5138
rect 152026 5057 152287 5097
rect 152026 5036 152047 5057
rect 151877 5020 152047 5036
rect 149908 4050 150268 4090
rect 149908 2940 149948 4050
rect 151877 3510 152047 3526
rect 151877 3408 151893 3510
rect 152026 3474 152047 3510
rect 152026 3434 152167 3474
rect 152026 3408 152047 3434
rect 151877 3392 152047 3408
rect 149902 2930 149954 2940
rect 149902 2722 149954 2730
rect 151877 1882 152047 1898
rect 151877 1780 151893 1882
rect 152026 1780 152047 1882
rect 151877 1764 152047 1780
rect 152007 678 152047 1764
rect 152127 678 152167 3434
rect 152247 678 152287 5057
rect 152367 678 152407 6699
rect 152500 6196 152540 7138
rect 152494 6186 152546 6196
rect 152494 5978 152546 5986
rect 152634 5870 152674 10786
rect 152500 5830 152674 5870
rect 152500 4568 152540 5830
rect 152494 4558 152546 4568
rect 152494 4350 152546 4358
rect 152820 4090 152860 10882
rect 154956 7178 154996 10978
rect 155092 7824 155132 11074
rect 155086 7814 155138 7824
rect 155086 7606 155138 7614
rect 154956 7138 155132 7178
rect 154469 6766 154639 6782
rect 154469 6664 154485 6766
rect 154618 6739 154639 6766
rect 154618 6699 154999 6739
rect 154618 6664 154639 6699
rect 154469 6648 154639 6664
rect 154469 5138 154639 5154
rect 154469 5036 154485 5138
rect 154618 5097 154639 5138
rect 154618 5057 154879 5097
rect 154618 5036 154639 5057
rect 154469 5020 154639 5036
rect 152500 4050 152860 4090
rect 152500 2940 152540 4050
rect 154469 3510 154639 3526
rect 154469 3408 154485 3510
rect 154618 3474 154639 3510
rect 154618 3434 154759 3474
rect 154618 3408 154639 3434
rect 154469 3392 154639 3408
rect 152494 2930 152546 2940
rect 152494 2722 152546 2730
rect 154469 1882 154639 1898
rect 154469 1780 154485 1882
rect 154618 1780 154639 1882
rect 154469 1764 154639 1780
rect 154599 678 154639 1764
rect 154719 678 154759 3434
rect 154839 678 154879 5057
rect 154959 678 154999 6699
rect 155092 6196 155132 7138
rect 155086 6186 155138 6196
rect 155086 5978 155138 5986
rect 155226 5870 155266 11170
rect 155092 5830 155266 5870
rect 155092 4568 155132 5830
rect 155086 4558 155138 4568
rect 155086 4350 155138 4358
rect 155412 4090 155452 11266
rect 157061 6766 157231 6782
rect 157061 6664 157077 6766
rect 157210 6739 157231 6766
rect 157210 6699 157591 6739
rect 157210 6664 157231 6699
rect 157061 6648 157231 6664
rect 157061 5138 157231 5154
rect 157061 5036 157077 5138
rect 157210 5097 157231 5138
rect 157210 5057 157471 5097
rect 157210 5036 157231 5057
rect 157061 5020 157231 5036
rect 155092 4050 155452 4090
rect 155092 2940 155132 4050
rect 157061 3510 157231 3526
rect 157061 3408 157077 3510
rect 157210 3474 157231 3510
rect 157210 3434 157351 3474
rect 157210 3408 157231 3434
rect 157061 3392 157231 3408
rect 155086 2930 155138 2940
rect 155086 2722 155138 2730
rect 157061 1882 157231 1898
rect 157061 1780 157077 1882
rect 157210 1780 157231 1882
rect 157061 1764 157231 1780
rect 157191 678 157231 1764
rect 157311 678 157351 3434
rect 157431 678 157471 5057
rect 157551 678 157591 6699
rect 130336 112 139084 152
<< via2 >>
rect 92448 8465 92775 8697
rect 103368 8465 103695 8697
rect 105264 8465 105591 8697
rect 111138 8465 111465 8697
rect 113274 8465 113601 8697
rect 114342 8465 114669 8697
rect 120750 8465 121077 8697
rect 125556 8465 125883 8697
rect 127158 8465 127485 8697
rect 128760 8465 129087 8697
rect 130362 8465 130689 8697
rect 131964 8465 132291 8697
rect 133566 8465 133893 8697
rect 135168 8465 135495 8697
rect 135997 8465 136169 8697
rect 137655 7426 137910 7660
rect 83084 4654 137146 4738
rect 137654 4638 137909 4872
rect 138108 4657 138215 6299
rect 83084 4379 137147 4463
rect 83162 4377 109062 4379
rect 138379 1342 138593 2481
rect 137068 1099 137185 1287
rect 129222 843 129549 1031
rect 132450 843 132777 1031
rect 133529 843 133856 1031
rect 134534 843 134861 1031
rect 135582 843 135909 1031
rect 140035 1563 141277 2485
rect 140035 1448 141277 1563
rect 140035 1340 141277 1448
rect 142647 5637 143849 6280
rect 142647 5420 143849 5637
rect 142647 4689 143849 5420
rect 145367 7003 146299 7851
rect 145367 6946 146299 7003
rect 145367 6713 146299 6946
<< metal3 >>
rect 92431 8697 92789 11254
rect 103111 9436 103469 11254
rect 103110 9426 103470 9436
rect 103110 9115 103123 9426
rect 103456 9378 103470 9426
rect 103456 9115 103709 9378
rect 103110 9100 103709 9115
rect 103111 9020 103709 9100
rect 92431 8465 92448 8697
rect 92775 8465 92789 8697
rect 92431 8444 92789 8465
rect 103351 8697 103709 9020
rect 103351 8465 103368 8697
rect 103695 8465 103709 8697
rect 103351 8444 103709 8465
rect 105247 8697 105605 11254
rect 105247 8465 105264 8697
rect 105591 8465 105605 8697
rect 105247 8444 105605 8465
rect 111121 9937 111479 11254
rect 111121 9633 111131 9937
rect 111469 9633 111479 9937
rect 111121 8697 111479 9633
rect 111121 8465 111138 8697
rect 111465 8465 111479 8697
rect 111121 8444 111479 8465
rect 113257 9453 113615 11254
rect 113257 9149 113265 9453
rect 113603 9149 113615 9453
rect 113257 8697 113615 9149
rect 113257 8465 113274 8697
rect 113601 8465 113615 8697
rect 113257 8444 113615 8465
rect 114325 8697 114683 11254
rect 114325 8465 114342 8697
rect 114669 8465 114683 8697
rect 114325 8444 114683 8465
rect 120733 8697 121091 11254
rect 120733 8465 120750 8697
rect 121077 8465 121091 8697
rect 120733 8444 121091 8465
rect 125539 8977 125897 11254
rect 125539 8685 125554 8977
rect 125882 8697 125897 8977
rect 125539 8465 125556 8685
rect 125883 8465 125897 8697
rect 125539 8453 125897 8465
rect 127141 8697 127499 11254
rect 127141 8465 127158 8697
rect 127485 8465 127499 8697
rect 127141 8444 127499 8465
rect 128743 8697 129101 11254
rect 128743 8465 128760 8697
rect 129087 8465 129101 8697
rect 128743 8444 129101 8465
rect 130345 8697 130703 11254
rect 130345 8465 130362 8697
rect 130689 8465 130703 8697
rect 130345 8444 130703 8465
rect 131947 8697 132305 11254
rect 131947 8465 131964 8697
rect 132291 8465 132305 8697
rect 131947 8444 132305 8465
rect 133549 8697 133907 11254
rect 133549 8465 133566 8697
rect 133893 8465 133907 8697
rect 133549 8444 133907 8465
rect 135151 8697 135509 11254
rect 135151 8465 135168 8697
rect 135495 8465 135509 8697
rect 135151 8444 135509 8465
rect 135980 8697 136219 11254
rect 142069 9922 142414 9933
rect 142069 9639 142084 9922
rect 142407 9639 142414 9922
rect 141505 9444 141850 9463
rect 141505 9155 141519 9444
rect 141839 9155 141850 9444
rect 135980 8465 135997 8697
rect 136169 8465 136219 8697
rect 135980 8444 136219 8465
rect 139415 8974 139760 8983
rect 139415 8685 139427 8974
rect 139747 8685 139760 8974
rect 138784 8446 139129 8461
rect 138784 8151 138802 8446
rect 139118 8151 139129 8446
rect 137642 7660 137920 7697
rect 137642 7426 137655 7660
rect 137910 7426 137920 7660
rect 137642 4872 137920 7426
rect 82876 4827 137654 4872
rect 82876 4653 83084 4827
rect 137147 4653 137654 4827
rect 82876 4638 137654 4653
rect 137909 4638 137920 4872
rect 138079 6299 138248 6321
rect 138079 4657 138108 6299
rect 138215 4657 138248 6299
rect 138079 4638 138248 4657
rect 82887 4464 137539 4480
rect 82887 4290 83084 4464
rect 137147 4290 137539 4464
rect 82887 4288 83162 4290
rect 109062 4288 137539 4290
rect 82887 4242 137539 4288
rect 137642 1493 137920 4638
rect 138358 2481 138622 2512
rect 138358 1342 138379 2481
rect 138593 1342 138622 2481
rect 138358 1310 138622 1342
rect 137060 1287 137194 1303
rect 137060 1099 137068 1287
rect 137185 1099 137194 1287
rect 137060 1092 137194 1099
rect 129205 1031 129567 1053
rect 129205 843 129222 1031
rect 129549 843 129567 1031
rect 129205 379 129567 843
rect 132433 1031 132795 1053
rect 132433 843 132450 1031
rect 132777 843 132795 1031
rect 129205 369 129584 379
rect 129205 19 129223 369
rect 129573 19 129584 369
rect 129205 0 129584 19
rect 132433 0 132795 843
rect 133512 1031 133874 1053
rect 133512 843 133529 1031
rect 133856 843 133874 1031
rect 133512 367 133874 843
rect 133512 12 133520 367
rect 133864 12 133874 367
rect 133512 1 133874 12
rect 134517 1031 134879 1053
rect 134517 843 134534 1031
rect 134861 843 134879 1031
rect 134517 363 134879 843
rect 135565 1031 135923 1053
rect 135565 843 135582 1031
rect 135909 843 135923 1031
rect 135565 803 135923 843
rect 135565 778 135927 803
rect 138784 778 139129 8151
rect 135565 447 139129 778
rect 139415 363 139760 8685
rect 140009 2485 141309 2513
rect 140009 1340 140035 2485
rect 141277 1340 141309 2485
rect 140009 1313 141309 1340
rect 141505 381 141850 9155
rect 142069 957 142414 9639
rect 145336 7851 146329 7886
rect 145336 6713 145367 7851
rect 146299 6713 146329 7851
rect 145336 6684 146329 6713
rect 142588 6280 143894 6323
rect 142588 4689 142647 6280
rect 143849 4689 143894 6280
rect 142588 4636 143894 4689
rect 142069 609 142086 957
rect 142404 609 142414 957
rect 142069 592 142414 609
rect 134517 1 139760 363
rect 141503 365 141850 381
rect 141503 17 141518 365
rect 141836 17 141850 365
rect 141503 0 141850 17
<< via3 >>
rect 103123 9115 103456 9426
rect 111131 9633 111469 9937
rect 113265 9149 113603 9453
rect 125554 8697 125882 8977
rect 125554 8685 125556 8697
rect 125556 8685 125882 8697
rect 142084 9639 142407 9922
rect 141519 9155 141839 9444
rect 139427 8685 139747 8974
rect 138802 8151 139118 8446
rect 83084 4738 137147 4827
rect 83084 4654 137146 4738
rect 137146 4654 137147 4738
rect 83084 4653 137147 4654
rect 138108 4657 138215 6299
rect 83084 4463 137147 4464
rect 83084 4379 137147 4463
rect 83084 4377 83162 4379
rect 83162 4377 109062 4379
rect 109062 4377 137147 4379
rect 83084 4290 137147 4377
rect 83162 4288 109062 4290
rect 138379 1342 138593 2481
rect 129223 19 129573 369
rect 133520 12 133864 367
rect 140035 1340 141277 2485
rect 145367 6713 146299 7851
rect 142647 4689 143849 6280
rect 142086 609 142404 957
rect 141518 17 141836 365
<< metal4 >>
rect 111113 9937 142416 9942
rect 111113 9633 111131 9937
rect 111469 9922 142416 9937
rect 111469 9639 142084 9922
rect 142407 9639 142416 9922
rect 111469 9633 142416 9639
rect 111113 9622 142416 9633
rect 113256 9453 141850 9462
rect 103110 9426 103470 9436
rect 103110 9115 103123 9426
rect 103456 9115 103470 9426
rect 113256 9149 113265 9453
rect 113603 9444 141850 9453
rect 113603 9155 141519 9444
rect 141839 9155 141850 9444
rect 113603 9149 141850 9155
rect 113256 9142 141850 9149
rect 103110 9100 103470 9115
rect 103147 8458 103467 9100
rect 125536 8977 139756 8992
rect 125536 8685 125554 8977
rect 125882 8974 139756 8977
rect 125882 8685 139427 8974
rect 139747 8685 139756 8974
rect 125536 8672 139756 8685
rect 103147 8446 139135 8458
rect 103147 8151 138802 8446
rect 139118 8151 139135 8446
rect 103147 8138 139135 8151
rect 138356 7851 157853 7883
rect 138356 6713 145367 7851
rect 146299 6713 157853 7851
rect 138356 6683 157853 6713
rect 82835 6299 157853 6320
rect 82835 4827 138108 6299
rect 82835 4653 83084 4827
rect 137147 4657 138108 4827
rect 138215 6280 157853 6299
rect 138215 4689 142647 6280
rect 143849 4689 157853 6280
rect 138215 4657 157853 4689
rect 137147 4653 157853 4657
rect 82835 4635 157853 4653
rect 82836 4464 157853 4484
rect 82836 4290 83084 4464
rect 137147 4290 157853 4464
rect 82836 4288 83162 4290
rect 109062 4288 157853 4290
rect 82836 2799 157853 4288
rect 138356 2485 157853 2511
rect 138356 2481 140035 2485
rect 138356 1342 138379 2481
rect 138593 1342 140035 2481
rect 138356 1340 140035 1342
rect 141277 1340 157853 2485
rect 138356 1311 157853 1340
rect 129205 957 142419 971
rect 129205 609 142086 957
rect 142404 609 142419 957
rect 129205 592 142419 609
rect 129205 369 129584 592
rect 141503 380 141850 381
rect 129205 19 129223 369
rect 129573 19 129584 369
rect 129205 0 129584 19
rect 133512 367 141850 380
rect 133512 12 133520 367
rect 133864 365 141850 367
rect 133864 17 141518 365
rect 141836 17 141850 365
rect 133864 12 141850 17
rect 133512 1 141850 12
rect 141503 0 141850 1
use bias_nstack  bias_nstack_0
array 0 101 -534 0 0 -3895
timestamp 1747745286
transform -1 0 86919 0 -1 1620
box 3258 -2860 3926 785
use bias_pstack  bias_pstack_0
array 0 101 534 0 0 -3895
timestamp 1747745073
transform 1 0 80966 0 -1 5026
box 1986 -3697 2714 338
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1746753973
transform -1 0 139896 0 -1 4714
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_1
timestamp 1746753973
transform -1 0 139896 0 -1 7970
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_14
timestamp 1746753973
transform -1 0 139896 0 -1 3086
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_18
timestamp 1746753973
transform -1 0 139896 0 -1 6342
box -66 -43 450 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1746753973
transform 1 0 139704 0 1 1458
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_1
timestamp 1746753973
transform 1 0 155256 0 1 1458
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_2
timestamp 1746753973
transform 1 0 152664 0 1 1458
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_3
timestamp 1746753973
transform 1 0 150072 0 1 1458
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_4
timestamp 1746753973
transform 1 0 147480 0 1 1458
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_5
timestamp 1746753973
transform 1 0 144888 0 1 1458
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_6
timestamp 1746753973
transform 1 0 142296 0 1 1458
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_7
timestamp 1746753973
transform 1 0 139704 0 1 4714
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_8
timestamp 1746753973
transform 1 0 139704 0 1 3086
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_9
timestamp 1746753973
transform 1 0 139704 0 1 6342
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_10
timestamp 1746753973
transform 1 0 142296 0 1 6342
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_11
timestamp 1746753973
transform 1 0 144888 0 1 6342
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_12
timestamp 1746753973
transform 1 0 147480 0 1 6342
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_13
timestamp 1746753973
transform 1 0 150072 0 1 6342
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_14
timestamp 1746753973
transform 1 0 152664 0 1 6342
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_15
timestamp 1746753973
transform 1 0 142296 0 1 4714
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_16
timestamp 1746753973
transform 1 0 155256 0 1 6342
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_17
timestamp 1746753973
transform 1 0 155256 0 1 4714
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_18
timestamp 1746753973
transform 1 0 155256 0 1 3086
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_19
timestamp 1746753973
transform 1 0 152664 0 1 3086
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_20
timestamp 1746753973
transform 1 0 150072 0 1 3086
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_21
timestamp 1746753973
transform 1 0 147480 0 1 3086
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_22
timestamp 1746753973
transform 1 0 144888 0 1 3086
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_23
timestamp 1746753973
transform 1 0 142296 0 1 3086
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_24
timestamp 1746753973
transform 1 0 144888 0 1 4714
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_25
timestamp 1746753973
transform 1 0 147480 0 1 4714
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_26
timestamp 1746753973
transform 1 0 150072 0 1 4714
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_27
timestamp 1746753973
transform 1 0 152664 0 1 4714
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1746753973
transform -1 0 144696 0 1 1458
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_1
timestamp 1746753973
transform -1 0 149880 0 1 4714
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_2
timestamp 1746753973
transform -1 0 149880 0 1 3086
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_3
timestamp 1746753973
transform -1 0 147288 0 1 1458
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_4
timestamp 1746753973
transform -1 0 144696 0 1 6342
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_5
timestamp 1746753973
transform -1 0 149880 0 1 6342
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_6
timestamp 1746753973
transform -1 0 144696 0 1 4714
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_7
timestamp 1746753973
transform -1 0 144696 0 1 3086
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_8
timestamp 1746753973
transform -1 0 142104 0 1 1458
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_9
timestamp 1746753973
transform -1 0 142104 0 1 4714
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_10
timestamp 1746753973
transform -1 0 142104 0 1 3086
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_11
timestamp 1746753973
transform -1 0 139512 0 1 1458
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_12
timestamp 1746753973
transform -1 0 142104 0 1 6342
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_13
timestamp 1746753973
transform -1 0 139512 0 1 6342
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_14
timestamp 1746753973
transform -1 0 139512 0 -1 3086
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_15
timestamp 1746753973
transform -1 0 139512 0 -1 4714
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_16
timestamp 1746753973
transform -1 0 139512 0 1 4714
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_17
timestamp 1746753973
transform -1 0 139512 0 1 3086
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_18
timestamp 1746753973
transform -1 0 139512 0 -1 6342
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_19
timestamp 1746753973
transform -1 0 139512 0 -1 7970
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_20
timestamp 1746753973
transform -1 0 149880 0 1 1458
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_21
timestamp 1746753973
transform -1 0 147288 0 1 3086
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_22
timestamp 1746753973
transform -1 0 147288 0 1 4714
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_23
timestamp 1746753973
transform -1 0 147288 0 1 6342
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_24
timestamp 1746753973
transform -1 0 155064 0 1 1458
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_25
timestamp 1746753973
transform -1 0 155064 0 1 6342
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_26
timestamp 1746753973
transform -1 0 155064 0 1 4714
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_27
timestamp 1746753973
transform -1 0 155064 0 1 3086
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_28
timestamp 1746753973
transform -1 0 152472 0 1 1458
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_29
timestamp 1746753973
transform -1 0 152472 0 1 6342
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_30
timestamp 1746753973
transform -1 0 152472 0 1 4714
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_31
timestamp 1746753973
transform -1 0 152472 0 1 3086
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1746753973
transform 1 0 139512 0 1 1458
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_1
timestamp 1746753973
transform 1 0 155064 0 1 1458
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_2
timestamp 1746753973
transform 1 0 152472 0 1 1458
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_3
timestamp 1746753973
transform 1 0 149880 0 1 1458
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_4
timestamp 1746753973
transform 1 0 147288 0 1 1458
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_5
timestamp 1746753973
transform 1 0 144696 0 1 1458
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_6
timestamp 1746753973
transform 1 0 142104 0 1 1458
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_7
timestamp 1746753973
transform 1 0 139512 0 1 4714
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_8
timestamp 1746753973
transform 1 0 139512 0 1 3086
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_9
timestamp 1746753973
transform 1 0 139512 0 1 6342
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_10
timestamp 1746753973
transform 1 0 142104 0 1 6342
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_11
timestamp 1746753973
transform 1 0 144696 0 1 6342
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_12
timestamp 1746753973
transform 1 0 147288 0 1 6342
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_13
timestamp 1746753973
transform 1 0 149880 0 1 6342
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_14
timestamp 1746753973
transform 1 0 152472 0 1 6342
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_15
timestamp 1746753973
transform 1 0 142104 0 1 4714
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_16
timestamp 1746753973
transform 1 0 155064 0 1 6342
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_17
timestamp 1746753973
transform 1 0 155064 0 1 4714
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_18
timestamp 1746753973
transform 1 0 155064 0 1 3086
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_19
timestamp 1746753973
transform 1 0 152472 0 1 3086
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_20
timestamp 1746753973
transform 1 0 149880 0 1 3086
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_21
timestamp 1746753973
transform 1 0 147288 0 1 3086
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_22
timestamp 1746753973
transform 1 0 144696 0 1 3086
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_23
timestamp 1746753973
transform 1 0 142104 0 1 3086
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_24
timestamp 1746753973
transform 1 0 144696 0 1 4714
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_25
timestamp 1746753973
transform 1 0 147288 0 1 4714
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_26
timestamp 1746753973
transform 1 0 149880 0 1 4714
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_27
timestamp 1746753973
transform 1 0 152472 0 1 4714
box -66 -43 258 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1746753973
transform -1 0 142488 0 -1 3086
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_1
timestamp 1746753973
transform -1 0 145080 0 -1 4714
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_2
timestamp 1746753973
transform -1 0 150264 0 -1 7970
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_3
timestamp 1746753973
transform -1 0 150264 0 -1 6342
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_4
timestamp 1746753973
transform -1 0 150264 0 -1 4714
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_5
timestamp 1746753973
transform -1 0 145080 0 -1 7970
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_6
timestamp 1746753973
transform -1 0 145080 0 -1 6342
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_7
timestamp 1746753973
transform -1 0 142488 0 -1 4714
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_8
timestamp 1746753973
transform -1 0 147672 0 -1 3086
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_9
timestamp 1746753973
transform -1 0 150264 0 -1 3086
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_10
timestamp 1746753973
transform -1 0 142488 0 -1 7970
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_11
timestamp 1746753973
transform -1 0 142488 0 -1 6342
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_12
timestamp 1746753973
transform -1 0 145080 0 -1 3086
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_13
timestamp 1746753973
transform -1 0 147672 0 -1 4714
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_14
timestamp 1746753973
transform -1 0 147672 0 -1 6342
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_15
timestamp 1746753973
transform -1 0 147672 0 -1 7970
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_16
timestamp 1746753973
transform -1 0 155448 0 -1 3086
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_17
timestamp 1746753973
transform -1 0 155448 0 -1 7970
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_18
timestamp 1746753973
transform -1 0 155448 0 -1 6342
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_19
timestamp 1746753973
transform -1 0 155448 0 -1 4714
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_20
timestamp 1746753973
transform -1 0 152856 0 -1 3086
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_21
timestamp 1746753973
transform -1 0 152856 0 -1 7970
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_22
timestamp 1746753973
transform -1 0 152856 0 -1 6342
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_23
timestamp 1746753973
transform -1 0 152856 0 -1 4714
box -66 -43 546 897
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
array 0 6 -2592 0 3 1628
timestamp 1746753973
transform -1 0 142008 0 1 1458
box -66 -43 2178 1671
<< labels >>
flabel metal4 157253 1311 157853 2511 0 FreeSans 3200 90 0 0 dvss
port 4 nsew
flabel metal4 157253 2799 157853 4484 0 FreeSans 3200 90 0 0 avss
port 2 nsew
flabel metal4 157253 4635 157853 6320 0 FreeSans 3200 90 0 0 avdd
port 1 nsew
flabel metal4 157253 6683 157853 7883 0 FreeSans 3200 90 0 0 dvdd
port 3 nsew
flabel metal3 92431 10225 92789 10465 0 FreeSans 1600 90 0 0 idac_src_1000
port 38 nsew
flabel metal3 111121 10225 111479 10465 0 FreeSans 1600 90 0 0 test_src_500
port 36 nsew
flabel metal3 113257 10225 113615 10465 0 FreeSans 1600 90 0 0 user_src_150
port 35 nsew
flabel metal3 114325 10225 114683 10465 0 FreeSans 1600 90 0 0 user_src_50
port 34 nsew
flabel metal3 120733 10225 121091 10465 0 FreeSans 1600 90 0 0 ov_src_600
port 33 nsew
flabel metal3 127141 10225 127499 10465 0 FreeSans 1600 90 0 0 instr2_src_100
port 31 nsew
flabel metal3 128743 10225 129101 10465 0 FreeSans 1600 90 0 0 instr1_src_100
port 30 nsew
flabel metal3 130345 10225 130703 10465 0 FreeSans 1600 90 0 0 hgbw2_src_100
port 29 nsew
flabel metal3 131947 10225 132305 10465 0 FreeSans 1600 90 0 0 hgbw1_src_100
port 28 nsew
flabel metal3 133549 10225 133907 10465 0 FreeSans 1600 90 0 0 lp2_src_100
port 27 nsew
flabel metal3 135151 10225 135509 10465 0 FreeSans 1600 90 0 0 lp1_src_100
port 8 nsew
flabel metal3 135980 10225 136219 10465 0 FreeSans 1600 90 0 0 lsxo_src_50
port 7 nsew
flabel metal2 157551 678 157591 1053 0 FreeSans 400 90 0 0 en_hsxo_bias
port 18 nsew
flabel metal2 157311 678 157351 1053 0 FreeSans 400 90 0 0 en_hsxo_trim_p
port 17 nsew
flabel metal2 157191 678 157231 1053 0 FreeSans 400 90 0 0 en_idac_bias
port 39 nsew
flabel metal2 154959 678 154999 1052 0 FreeSans 400 90 0 0 en_user2_bias
port 40 nsew
flabel metal2 154839 678 154879 1052 0 FreeSans 400 90 0 0 en_user1_bias
port 41 nsew
flabel metal2 154719 678 154759 1052 0 FreeSans 400 90 0 0 en_user2_trim_p
port 42 nsew
flabel metal2 154599 678 154639 1052 0 FreeSans 400 90 0 0 en_src_test
port 43 nsew
flabel metal2 152367 678 152407 1052 0 FreeSans 400 90 0 0 en_comp_bias
port 44 nsew
flabel metal2 152247 678 152287 1052 0 FreeSans 400 90 0 0 en_instr2_trim_p
port 45 nsew
flabel metal2 152127 678 152167 1052 0 FreeSans 400 90 0 0 en_comp_trim_p
port 46 nsew
flabel metal2 152007 678 152047 1052 0 FreeSans 400 90 0 0 en_ov_bias
port 47 nsew
flabel metal2 149775 678 149815 1052 0 FreeSans 400 90 0 0 en_instr1_bias
port 48 nsew
flabel metal2 149655 678 149695 1052 0 FreeSans 400 90 0 0 en_hgbw2_trim_p
port 49 nsew
flabel metal2 149535 678 149575 1052 0 FreeSans 400 90 0 0 en_instr1_trim_p
port 50 nsew
flabel metal2 149415 678 149455 1052 0 FreeSans 400 90 0 0 en_instr2_bias
port 51 nsew
flabel metal2 147183 678 147223 1051 0 FreeSans 400 90 0 0 en_hgbw1_bias
port 52 nsew
flabel metal2 147063 678 147103 1051 0 FreeSans 400 90 0 0 en_lp2_trim_p
port 53 nsew
flabel metal2 146943 678 146983 1051 0 FreeSans 400 90 0 0 en_hgbw1_trim_p
port 54 nsew
flabel metal2 146823 678 146863 1051 0 FreeSans 400 90 0 0 en_hgbw2_bias
port 55 nsew
flabel metal2 144591 678 144631 1053 0 FreeSans 400 90 0 0 en_lp1_bias
port 22 nsew
flabel metal2 144471 678 144511 1053 0 FreeSans 400 90 0 0 en_lsxo_bias
port 23 nsew
flabel metal2 144351 678 144391 1053 0 FreeSans 400 90 0 0 en_lp1_trim_p
port 21 nsew
flabel metal2 144231 678 144271 1053 0 FreeSans 400 90 0 0 en_lp2_bias
port 20 nsew
flabel metal2 141999 678 142039 1053 0 FreeSans 400 90 0 0 en_hsxo_trim_n
port 25 nsew
flabel metal2 141879 678 141919 1053 0 FreeSans 400 90 0 0 en_comp_trim_n
port 24 nsew
flabel metal2 141763 678 141803 1053 0 FreeSans 400 90 0 0 en_user2_trim_n
port 16 nsew
flabel metal2 141639 678 141679 1078 0 FreeSans 400 90 0 0 en_snk_test
port 26 nsew
flabel metal2 157431 678 157471 1053 0 FreeSans 400 90 0 0 en_brnout_bias
port 19 nsew
flabel metal4 82835 4635 83068 6320 0 FreeSans 1600 90 0 0 avdd
port 1 nsew
flabel metal3 105247 10225 105605 10465 0 FreeSans 1600 90 0 0 brnout_src_200
port 56 nsew
flabel metal4 82836 2799 83069 4484 0 FreeSans 1600 90 0 0 avss
port 2 nsew
flabel metal3 125539 10225 125897 10465 0 FreeSans 1600 90 0 0 comp_src_400
port 32 nsew
flabel metal3 132433 0 132795 291 0 FreeSans 1600 90 0 0 bandgap_snk_250
port 58 nsew
flabel metal3 103111 10225 103469 10465 0 FreeSans 1600 90 0 0 hsxo_src_100
port 37 nsew
<< properties >>
string MASKHINTS_HVI 139065 1215 157825 1485 139060 7965 157820 8235 139090 1250 139735 8190 157430 1260 157835 8190
<< end >>
