magic
tech sky130A
magscale 1 2
timestamp 1719795003
<< viali >>
rect 1092 1950 1160 2854
<< metal1 >>
rect 435 7250 5527 7371
rect 856 4999 1044 5067
rect 852 3371 1040 3439
rect 1078 3438 1162 3440
rect 1078 2854 1174 3438
rect 1078 1950 1092 2854
rect 1160 1950 1174 2854
rect 1078 1746 1174 1950
<< metal2 >>
rect 47877 7213 48035 7273
<< via2 >>
rect 7681 34828 47745 34890
rect 7699 26652 47763 26714
rect 1005 25695 47470 25757
rect 1553 17526 41617 17588
rect 1028 16343 41092 16405
rect 1005 8161 47469 8223
rect 45880 7213 47877 7273
rect 45884 -946 48005 -888
<< metal3 >>
rect 49073 34950 49433 35112
rect 7638 34890 49433 34950
rect 7638 34828 7681 34890
rect 47745 34828 49433 34890
rect 7638 34758 49433 34828
rect 7648 26773 48043 26812
rect 7648 26714 47837 26773
rect 7648 26652 7699 26714
rect 47763 26652 47837 26714
rect 7648 26576 47837 26652
rect 47807 25858 47837 26576
rect 951 25757 47837 25858
rect 951 25695 1005 25757
rect 47470 25695 47837 25757
rect 951 25639 47837 25695
rect 47999 25639 48043 26773
rect 951 25599 48043 25639
rect 951 25597 48033 25599
rect 49073 17659 49433 34758
rect 1478 17588 49433 17659
rect 1478 17526 1553 17588
rect 41617 17526 49433 17588
rect 1478 17464 49433 17526
rect 47867 16464 49433 17464
rect 978 16405 49433 16464
rect 978 16343 1028 16405
rect 41092 16343 49433 16405
rect 978 16269 49433 16343
rect 960 8267 48113 8312
rect 960 8223 47902 8267
rect 960 8161 1005 8223
rect 47469 8161 47902 8223
rect 960 8087 47902 8161
rect 47877 7363 47902 8087
rect 45838 7273 47902 7363
rect 45838 7213 45880 7273
rect 47877 7213 47902 7273
rect 45838 7154 47902 7213
rect 48078 7154 48113 8267
rect 45838 7127 48113 7154
rect 49073 -824 49433 16269
rect 45847 -888 49433 -824
rect 45847 -946 45884 -888
rect 48005 -946 49433 -888
rect 45847 -1007 49433 -946
rect 4254 -1161 19726 -1041
rect 49073 -1043 49433 -1007
rect 49553 26768 49913 35112
rect 49553 25637 49590 26768
rect 49868 25637 49913 26768
rect 49553 8277 49913 25637
rect 49553 7154 49577 8277
rect 49886 7154 49913 8277
rect 49553 -1043 49913 7154
<< via3 >>
rect 47837 25639 47999 26773
rect 47902 7154 48078 8267
rect 49590 25637 49868 26768
rect 49577 7154 49886 8277
<< metal4 >>
rect 47801 26773 49911 26814
rect 47801 25639 47837 26773
rect 47999 26768 49911 26773
rect 47999 25639 49590 26768
rect 47801 25637 49590 25639
rect 49868 25637 49911 26768
rect 47801 25601 49911 25637
rect 47875 8277 49917 8310
rect 47875 8267 49577 8277
rect 47875 7154 47902 8267
rect 48078 7154 49577 8267
rect 49886 7154 49917 8277
rect 47875 7123 49917 7154
use bias_generator_fe  bias_generator_fe_0
timestamp 1719596014
transform 1 0 -35 0 1 -1186
box 1072 0 45976 8863
use bias_generator_idac_be  bias_generator_idac_be_0
timestamp 1719794226
transform 1 0 -89608 0 1 9596
box 88136 -10736 138547 25480
<< end >>
