magic
tech sky130A
magscale 1 2
timestamp 1747752771
<< viali >>
rect 1082 218 1148 1710
<< metal1 >>
rect 435 7250 5527 7371
rect 856 4999 1685 5067
rect 1078 3439 1162 3440
rect 852 3371 1685 3439
rect 1037 1743 1685 1811
rect 1052 1710 1176 1743
rect 1052 218 1082 1710
rect 1148 218 1176 1710
rect 1052 183 1176 218
rect 1037 115 1685 183
<< metal2 >>
rect 142 34487 182 34862
rect 262 34487 302 34862
rect 382 34487 422 34862
rect 502 34487 542 34862
rect 2734 34487 2774 34862
rect 2854 34487 2894 34862
rect 2970 34487 3010 34862
rect 3094 34462 3134 34862
rect 48508 27061 49914 27080
rect 48508 25352 48529 27061
rect 48833 25352 49574 27061
rect 48508 25346 49574 25352
rect 49888 25346 49914 27061
rect 48508 25327 49914 25346
rect 47968 10123 48017 10357
rect 48511 8554 49913 8581
rect 48511 8550 49576 8554
rect 47877 6943 48035 7003
rect 48511 6890 48546 8550
rect 48816 6890 49576 8550
rect 48511 6880 49576 6890
rect 49888 6880 49913 8554
rect 48511 6857 49913 6880
<< via2 >>
rect 7681 34578 47745 34640
rect 7699 26922 47763 26984
rect 1005 25425 47470 25487
rect 48529 25352 48833 27061
rect 49574 25346 49888 27061
rect 1553 17776 41617 17838
rect 1028 16093 41092 16155
rect 1005 8431 47469 8493
rect 45880 6943 47877 7003
rect 48546 6890 48816 8550
rect 49576 6880 49888 8554
rect 45884 -696 48005 -638
<< metal3 >>
rect 49073 34700 49433 35112
rect 7638 34640 49433 34700
rect 7638 34578 7681 34640
rect 47745 34578 49433 34640
rect 7638 34508 49433 34578
rect 0 34198 246 34232
rect 0 33050 30 34198
rect 220 33050 246 34198
rect 0 33026 246 33050
rect -1071 32721 -931 32804
rect -1071 31067 -1060 32721
rect -944 31067 -931 32721
rect -1071 27624 -931 31067
rect -1170 27484 -931 27624
rect -790 30886 -650 32768
rect -790 29232 -781 30886
rect -665 29232 -650 30886
rect -1170 21346 -1030 27484
rect -790 27306 -650 29232
rect -1170 19692 -1158 21346
rect -1042 19692 -1030 21346
rect -1170 14236 -1030 19692
rect -1170 12582 -1160 14236
rect -1044 12582 -1030 14236
rect -1170 7109 -1030 12582
rect -970 27166 -650 27306
rect -970 23181 -830 27166
rect -352 27080 -212 28868
rect -970 21527 -959 23181
rect -843 21527 -830 23181
rect -970 12398 -830 21527
rect -970 10744 -957 12398
rect -841 10744 -830 12398
rect -970 7359 -830 10744
rect -770 26940 -212 27080
rect -770 7594 -630 26940
rect 48 26880 188 33026
rect -570 26740 188 26880
rect 336 28858 482 28860
rect 336 28836 650 28858
rect 336 27678 360 28836
rect 624 27678 650 28836
rect 336 27658 650 27678
rect -570 19396 -430 26740
rect 336 26645 482 27658
rect 7648 27061 48859 27082
rect 7648 26984 48529 27061
rect 7648 26922 7699 26984
rect 47763 26922 48529 26984
rect 7648 26846 48529 26922
rect -337 26499 482 26645
rect -337 24701 -191 26499
rect 47807 25588 48529 26846
rect 951 25487 48529 25588
rect 951 25425 1005 25487
rect 47470 25425 48529 25487
rect 951 25352 48529 25425
rect 48833 25352 48859 27061
rect 951 25327 48859 25352
rect -337 24692 9 24701
rect -337 24562 -164 24692
rect -2 24562 9 24692
rect -337 24555 9 24562
rect -570 19136 8 19396
rect -570 18494 -430 19136
rect -278 18494 8 19136
rect -570 18184 8 18494
rect -570 15748 -430 18184
rect 49073 17909 49433 34508
rect 1478 17838 49433 17909
rect 1478 17776 1553 17838
rect 41617 17776 49433 17838
rect 1478 17714 49433 17776
rect 47867 16214 49433 17714
rect 978 16155 49433 16214
rect 978 16093 1028 16155
rect 41092 16093 49433 16155
rect 978 16019 49433 16093
rect -570 15452 12 15748
rect -570 14810 -430 15452
rect -276 14810 12 15452
rect -570 14536 12 14810
rect -570 7794 -430 14536
rect -342 9340 8 9352
rect -342 9222 -162 9340
rect -4 9222 8 9340
rect -342 9208 8 9222
rect -342 8014 -198 9208
rect 960 8550 48855 8582
rect 960 8493 48546 8550
rect 960 8431 1005 8493
rect 47469 8431 48546 8493
rect 960 8357 48546 8431
rect -342 7870 2058 8014
rect -570 7654 1690 7794
rect -770 7454 1290 7594
rect -970 7219 937 7359
rect -1170 6969 688 7109
rect 548 2866 688 6969
rect 548 1212 555 2866
rect 669 1212 688 2866
rect 548 1123 688 1212
rect 797 4702 937 7219
rect 1150 6316 1290 7454
rect 1116 6296 1370 6316
rect 1116 4936 1132 6296
rect 1344 4936 1370 6296
rect 1116 4920 1370 4936
rect 797 3047 809 4702
rect 924 3047 937 4702
rect 797 1138 937 3047
rect 1550 296 1690 7654
rect 1914 6318 2058 7870
rect 47877 7093 48546 8357
rect 45838 7003 48546 7093
rect 45838 6943 45880 7003
rect 47877 6943 48546 7003
rect 45838 6890 48546 6943
rect 48816 6890 48855 8550
rect 45838 6857 48855 6890
rect 1914 6272 2216 6318
rect 1914 4950 1948 6272
rect 2186 4950 2216 6272
rect 1914 4918 2216 4950
rect 49073 -574 49433 16019
rect 45847 -638 49433 -574
rect 45847 -696 45884 -638
rect 48005 -696 49433 -638
rect 45847 -757 49433 -696
rect 4254 -1161 19726 -1041
rect 49073 -1043 49433 -757
rect 49553 27061 49913 35112
rect 49553 25346 49574 27061
rect 49888 25346 49913 27061
rect 49553 8554 49913 25346
rect 49553 6880 49576 8554
rect 49888 6880 49913 8554
rect 49553 -1043 49913 6880
<< via3 >>
rect 30 33050 220 34198
rect -1060 31067 -944 32721
rect -781 29232 -665 30886
rect -1158 19692 -1042 21346
rect -1160 12582 -1044 14236
rect -959 21527 -843 23181
rect -957 10744 -841 12398
rect 360 27678 624 28836
rect -164 24562 -2 24692
rect -162 9222 -4 9340
rect 555 1212 669 2866
rect 1132 4936 1344 6296
rect 809 3047 924 4702
rect 1948 4950 2186 6272
<< metal4 >>
rect -984 23181 -169 23196
rect -984 21527 -959 23181
rect -843 21527 -169 23181
rect -984 21511 -169 21527
rect -1182 21346 -163 21360
rect -1182 19692 -1158 21346
rect -1042 19692 -163 21346
rect -1182 19675 -163 19692
rect -1186 14236 -167 14254
rect -1186 12582 -1160 14236
rect -1044 12582 -167 14236
rect -1186 12569 -167 12582
rect -976 12398 -167 12418
rect -976 10744 -957 12398
rect -841 10744 -167 12398
rect -976 10733 -167 10744
rect 1063 6296 1663 6318
rect 1063 4936 1132 6296
rect 1344 4936 1663 6296
rect 1063 4918 1663 4936
rect 778 4702 1663 4716
rect 778 3047 809 4702
rect 924 3047 1663 4702
rect 778 3031 1663 3047
rect 544 2866 1663 2880
rect 544 1212 555 2866
rect 669 1212 1663 2866
rect 544 1195 1663 1212
rect 1063 -564 1663 996
use bias_generator_fe  bias_generator_fe_0
timestamp 1747752771
transform 1 0 -35 0 1 -1186
box 1072 0 46056 8863
use bias_generator_idac_be  bias_generator_idac_be_0
timestamp 1747752771
transform 1 0 -89608 0 1 9596
box 88536 -10736 139522 25480
<< labels >>
flabel metal1 1037 3371 1437 3439 0 FreeSans 480 0 0 0 ena
port 53 nsew
flabel metal1 1037 4999 1437 5067 0 FreeSans 480 0 0 0 ref_sel_vbg
port 52 nsew
flabel metal1 435 7250 754 7371 0 FreeSans 640 0 0 0 vbg
port 54 nsew
flabel metal4 1063 -564 1547 996 0 FreeSans 3200 90 0 0 dvss
port 50 nsew
flabel metal4 1063 1195 1663 2880 0 FreeSans 3200 90 0 0 avss
port 12 nsew
flabel metal4 1063 3031 1663 4716 0 FreeSans 3200 90 0 0 avdd
port 59 nsew
flabel metal4 s 1063 4918 1663 6318 0 FreeSans 3200 90 0 0 dvdd
port 58 n
flabel metal3 49073 -1043 49433 -118 0 FreeSans 1600 90 0 0 snk_out
port 60 nsew
flabel metal3 49553 -1043 49913 -114 0 FreeSans 1600 90 0 0 src_out
port 61 nsew
flabel metal2 142 34487 182 34862 0 FreeSans 400 270 0 0 din[0]
port 22 nsew
flabel metal2 262 34487 302 34862 0 FreeSans 400 270 0 0 din[1]
port 23 nsew
flabel metal2 382 34487 422 34862 0 FreeSans 400 270 0 0 din[2]
port 21 nsew
flabel metal2 502 34487 542 34862 0 FreeSans 400 270 0 0 din[3]
port 20 nsew
flabel metal2 2734 34487 2774 34862 0 FreeSans 400 270 0 0 din[4]
port 25 nsew
flabel metal2 2854 34487 2894 34862 0 FreeSans 400 270 0 0 din[5]
port 24 nsew
flabel metal2 2970 34487 3010 34862 0 FreeSans 400 270 0 0 din[6]
port 16 nsew
flabel metal2 3094 34462 3134 34862 0 FreeSans 400 270 0 0 din[7]
port 26 nsew
flabel metal3 4254 -1161 4658 -1041 0 FreeSans 1120 0 0 0 ref_in
port 62 nsew
<< end >>
