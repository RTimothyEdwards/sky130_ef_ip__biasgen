magic
tech sky130A
magscale 1 2
timestamp 1716925149
<< pwell >>
rect -5679 -3582 5679 3582
<< psubdiff >>
rect -5643 3512 -5547 3546
rect 5547 3512 5643 3546
rect -5643 3450 -5609 3512
rect 5609 3450 5643 3512
rect -5643 -3512 -5609 -3450
rect 5609 -3512 5643 -3450
rect -5643 -3546 -5547 -3512
rect 5547 -3546 5643 -3512
<< psubdiffcont >>
rect -5547 3512 5547 3546
rect -5643 -3450 -5609 3450
rect 5609 -3450 5643 3450
rect -5547 -3546 5547 -3512
<< xpolycontact >>
rect -5513 2984 -5443 3416
rect -5513 -3416 -5443 -2984
rect -5347 2984 -5277 3416
rect -5347 -3416 -5277 -2984
rect -5181 2984 -5111 3416
rect -5181 -3416 -5111 -2984
rect -5015 2984 -4945 3416
rect -5015 -3416 -4945 -2984
rect -4849 2984 -4779 3416
rect -4849 -3416 -4779 -2984
rect -4683 2984 -4613 3416
rect -4683 -3416 -4613 -2984
rect -4517 2984 -4447 3416
rect -4517 -3416 -4447 -2984
rect -4351 2984 -4281 3416
rect -4351 -3416 -4281 -2984
rect -4185 2984 -4115 3416
rect -4185 -3416 -4115 -2984
rect -4019 2984 -3949 3416
rect -4019 -3416 -3949 -2984
rect -3853 2984 -3783 3416
rect -3853 -3416 -3783 -2984
rect -3687 2984 -3617 3416
rect -3687 -3416 -3617 -2984
rect -3521 2984 -3451 3416
rect -3521 -3416 -3451 -2984
rect -3355 2984 -3285 3416
rect -3355 -3416 -3285 -2984
rect -3189 2984 -3119 3416
rect -3189 -3416 -3119 -2984
rect -3023 2984 -2953 3416
rect -3023 -3416 -2953 -2984
rect -2857 2984 -2787 3416
rect -2857 -3416 -2787 -2984
rect -2691 2984 -2621 3416
rect -2691 -3416 -2621 -2984
rect -2525 2984 -2455 3416
rect -2525 -3416 -2455 -2984
rect -2359 2984 -2289 3416
rect -2359 -3416 -2289 -2984
rect -2193 2984 -2123 3416
rect -2193 -3416 -2123 -2984
rect -2027 2984 -1957 3416
rect -2027 -3416 -1957 -2984
rect -1861 2984 -1791 3416
rect -1861 -3416 -1791 -2984
rect -1695 2984 -1625 3416
rect -1695 -3416 -1625 -2984
rect -1529 2984 -1459 3416
rect -1529 -3416 -1459 -2984
rect -1363 2984 -1293 3416
rect -1363 -3416 -1293 -2984
rect -1197 2984 -1127 3416
rect -1197 -3416 -1127 -2984
rect -1031 2984 -961 3416
rect -1031 -3416 -961 -2984
rect -865 2984 -795 3416
rect -865 -3416 -795 -2984
rect -699 2984 -629 3416
rect -699 -3416 -629 -2984
rect -533 2984 -463 3416
rect -533 -3416 -463 -2984
rect -367 2984 -297 3416
rect -367 -3416 -297 -2984
rect -201 2984 -131 3416
rect -201 -3416 -131 -2984
rect -35 2984 35 3416
rect -35 -3416 35 -2984
rect 131 2984 201 3416
rect 131 -3416 201 -2984
rect 297 2984 367 3416
rect 297 -3416 367 -2984
rect 463 2984 533 3416
rect 463 -3416 533 -2984
rect 629 2984 699 3416
rect 629 -3416 699 -2984
rect 795 2984 865 3416
rect 795 -3416 865 -2984
rect 961 2984 1031 3416
rect 961 -3416 1031 -2984
rect 1127 2984 1197 3416
rect 1127 -3416 1197 -2984
rect 1293 2984 1363 3416
rect 1293 -3416 1363 -2984
rect 1459 2984 1529 3416
rect 1459 -3416 1529 -2984
rect 1625 2984 1695 3416
rect 1625 -3416 1695 -2984
rect 1791 2984 1861 3416
rect 1791 -3416 1861 -2984
rect 1957 2984 2027 3416
rect 1957 -3416 2027 -2984
rect 2123 2984 2193 3416
rect 2123 -3416 2193 -2984
rect 2289 2984 2359 3416
rect 2289 -3416 2359 -2984
rect 2455 2984 2525 3416
rect 2455 -3416 2525 -2984
rect 2621 2984 2691 3416
rect 2621 -3416 2691 -2984
rect 2787 2984 2857 3416
rect 2787 -3416 2857 -2984
rect 2953 2984 3023 3416
rect 2953 -3416 3023 -2984
rect 3119 2984 3189 3416
rect 3119 -3416 3189 -2984
rect 3285 2984 3355 3416
rect 3285 -3416 3355 -2984
rect 3451 2984 3521 3416
rect 3451 -3416 3521 -2984
rect 3617 2984 3687 3416
rect 3617 -3416 3687 -2984
rect 3783 2984 3853 3416
rect 3783 -3416 3853 -2984
rect 3949 2984 4019 3416
rect 3949 -3416 4019 -2984
rect 4115 2984 4185 3416
rect 4115 -3416 4185 -2984
rect 4281 2984 4351 3416
rect 4281 -3416 4351 -2984
rect 4447 2984 4517 3416
rect 4447 -3416 4517 -2984
rect 4613 2984 4683 3416
rect 4613 -3416 4683 -2984
rect 4779 2984 4849 3416
rect 4779 -3416 4849 -2984
rect 4945 2984 5015 3416
rect 4945 -3416 5015 -2984
rect 5111 2984 5181 3416
rect 5111 -3416 5181 -2984
rect 5277 2984 5347 3416
rect 5277 -3416 5347 -2984
rect 5443 2984 5513 3416
rect 5443 -3416 5513 -2984
<< ppolyres >>
rect -5513 -2984 -5443 2984
rect -5347 -2984 -5277 2984
rect -5181 -2984 -5111 2984
rect -5015 -2984 -4945 2984
rect -4849 -2984 -4779 2984
rect -4683 -2984 -4613 2984
rect -4517 -2984 -4447 2984
rect -4351 -2984 -4281 2984
rect -4185 -2984 -4115 2984
rect -4019 -2984 -3949 2984
rect -3853 -2984 -3783 2984
rect -3687 -2984 -3617 2984
rect -3521 -2984 -3451 2984
rect -3355 -2984 -3285 2984
rect -3189 -2984 -3119 2984
rect -3023 -2984 -2953 2984
rect -2857 -2984 -2787 2984
rect -2691 -2984 -2621 2984
rect -2525 -2984 -2455 2984
rect -2359 -2984 -2289 2984
rect -2193 -2984 -2123 2984
rect -2027 -2984 -1957 2984
rect -1861 -2984 -1791 2984
rect -1695 -2984 -1625 2984
rect -1529 -2984 -1459 2984
rect -1363 -2984 -1293 2984
rect -1197 -2984 -1127 2984
rect -1031 -2984 -961 2984
rect -865 -2984 -795 2984
rect -699 -2984 -629 2984
rect -533 -2984 -463 2984
rect -367 -2984 -297 2984
rect -201 -2984 -131 2984
rect -35 -2984 35 2984
rect 131 -2984 201 2984
rect 297 -2984 367 2984
rect 463 -2984 533 2984
rect 629 -2984 699 2984
rect 795 -2984 865 2984
rect 961 -2984 1031 2984
rect 1127 -2984 1197 2984
rect 1293 -2984 1363 2984
rect 1459 -2984 1529 2984
rect 1625 -2984 1695 2984
rect 1791 -2984 1861 2984
rect 1957 -2984 2027 2984
rect 2123 -2984 2193 2984
rect 2289 -2984 2359 2984
rect 2455 -2984 2525 2984
rect 2621 -2984 2691 2984
rect 2787 -2984 2857 2984
rect 2953 -2984 3023 2984
rect 3119 -2984 3189 2984
rect 3285 -2984 3355 2984
rect 3451 -2984 3521 2984
rect 3617 -2984 3687 2984
rect 3783 -2984 3853 2984
rect 3949 -2984 4019 2984
rect 4115 -2984 4185 2984
rect 4281 -2984 4351 2984
rect 4447 -2984 4517 2984
rect 4613 -2984 4683 2984
rect 4779 -2984 4849 2984
rect 4945 -2984 5015 2984
rect 5111 -2984 5181 2984
rect 5277 -2984 5347 2984
rect 5443 -2984 5513 2984
<< locali >>
rect -5643 3450 -5609 3546
rect 5609 3450 5643 3546
rect -5643 -3546 -5609 -3450
rect 5609 -3546 5643 -3450
<< viali >>
rect -5609 3512 -5547 3546
rect -5547 3512 5547 3546
rect 5547 3512 5609 3546
rect -5497 3001 -5459 3398
rect -5331 3001 -5293 3398
rect -5165 3001 -5127 3398
rect -4999 3001 -4961 3398
rect -4833 3001 -4795 3398
rect -4667 3001 -4629 3398
rect -4501 3001 -4463 3398
rect -4335 3001 -4297 3398
rect -4169 3001 -4131 3398
rect -4003 3001 -3965 3398
rect -3837 3001 -3799 3398
rect -3671 3001 -3633 3398
rect -3505 3001 -3467 3398
rect -3339 3001 -3301 3398
rect -3173 3001 -3135 3398
rect -3007 3001 -2969 3398
rect -2841 3001 -2803 3398
rect -2675 3001 -2637 3398
rect -2509 3001 -2471 3398
rect -2343 3001 -2305 3398
rect -2177 3001 -2139 3398
rect -2011 3001 -1973 3398
rect -1845 3001 -1807 3398
rect -1679 3001 -1641 3398
rect -1513 3001 -1475 3398
rect -1347 3001 -1309 3398
rect -1181 3001 -1143 3398
rect -1015 3001 -977 3398
rect -849 3001 -811 3398
rect -683 3001 -645 3398
rect -517 3001 -479 3398
rect -351 3001 -313 3398
rect -185 3001 -147 3398
rect -19 3001 19 3398
rect 147 3001 185 3398
rect 313 3001 351 3398
rect 479 3001 517 3398
rect 645 3001 683 3398
rect 811 3001 849 3398
rect 977 3001 1015 3398
rect 1143 3001 1181 3398
rect 1309 3001 1347 3398
rect 1475 3001 1513 3398
rect 1641 3001 1679 3398
rect 1807 3001 1845 3398
rect 1973 3001 2011 3398
rect 2139 3001 2177 3398
rect 2305 3001 2343 3398
rect 2471 3001 2509 3398
rect 2637 3001 2675 3398
rect 2803 3001 2841 3398
rect 2969 3001 3007 3398
rect 3135 3001 3173 3398
rect 3301 3001 3339 3398
rect 3467 3001 3505 3398
rect 3633 3001 3671 3398
rect 3799 3001 3837 3398
rect 3965 3001 4003 3398
rect 4131 3001 4169 3398
rect 4297 3001 4335 3398
rect 4463 3001 4501 3398
rect 4629 3001 4667 3398
rect 4795 3001 4833 3398
rect 4961 3001 4999 3398
rect 5127 3001 5165 3398
rect 5293 3001 5331 3398
rect 5459 3001 5497 3398
rect -5643 -2810 -5609 2810
rect 5609 -2810 5643 2810
rect -5497 -3398 -5459 -3001
rect -5331 -3398 -5293 -3001
rect -5165 -3398 -5127 -3001
rect -4999 -3398 -4961 -3001
rect -4833 -3398 -4795 -3001
rect -4667 -3398 -4629 -3001
rect -4501 -3398 -4463 -3001
rect -4335 -3398 -4297 -3001
rect -4169 -3398 -4131 -3001
rect -4003 -3398 -3965 -3001
rect -3837 -3398 -3799 -3001
rect -3671 -3398 -3633 -3001
rect -3505 -3398 -3467 -3001
rect -3339 -3398 -3301 -3001
rect -3173 -3398 -3135 -3001
rect -3007 -3398 -2969 -3001
rect -2841 -3398 -2803 -3001
rect -2675 -3398 -2637 -3001
rect -2509 -3398 -2471 -3001
rect -2343 -3398 -2305 -3001
rect -2177 -3398 -2139 -3001
rect -2011 -3398 -1973 -3001
rect -1845 -3398 -1807 -3001
rect -1679 -3398 -1641 -3001
rect -1513 -3398 -1475 -3001
rect -1347 -3398 -1309 -3001
rect -1181 -3398 -1143 -3001
rect -1015 -3398 -977 -3001
rect -849 -3398 -811 -3001
rect -683 -3398 -645 -3001
rect -517 -3398 -479 -3001
rect -351 -3398 -313 -3001
rect -185 -3398 -147 -3001
rect -19 -3398 19 -3001
rect 147 -3398 185 -3001
rect 313 -3398 351 -3001
rect 479 -3398 517 -3001
rect 645 -3398 683 -3001
rect 811 -3398 849 -3001
rect 977 -3398 1015 -3001
rect 1143 -3398 1181 -3001
rect 1309 -3398 1347 -3001
rect 1475 -3398 1513 -3001
rect 1641 -3398 1679 -3001
rect 1807 -3398 1845 -3001
rect 1973 -3398 2011 -3001
rect 2139 -3398 2177 -3001
rect 2305 -3398 2343 -3001
rect 2471 -3398 2509 -3001
rect 2637 -3398 2675 -3001
rect 2803 -3398 2841 -3001
rect 2969 -3398 3007 -3001
rect 3135 -3398 3173 -3001
rect 3301 -3398 3339 -3001
rect 3467 -3398 3505 -3001
rect 3633 -3398 3671 -3001
rect 3799 -3398 3837 -3001
rect 3965 -3398 4003 -3001
rect 4131 -3398 4169 -3001
rect 4297 -3398 4335 -3001
rect 4463 -3398 4501 -3001
rect 4629 -3398 4667 -3001
rect 4795 -3398 4833 -3001
rect 4961 -3398 4999 -3001
rect 5127 -3398 5165 -3001
rect 5293 -3398 5331 -3001
rect 5459 -3398 5497 -3001
rect -5609 -3546 -5547 -3512
rect -5547 -3546 5547 -3512
rect 5547 -3546 5609 -3512
<< metal1 >>
rect -5621 3546 5621 3552
rect -5621 3512 -5609 3546
rect 5609 3512 5621 3546
rect -5621 3506 5621 3512
rect -5503 3398 -5453 3410
rect -5503 3001 -5497 3398
rect -5459 3001 -5453 3398
rect -5503 2989 -5453 3001
rect -5337 3398 -5287 3410
rect -5337 3001 -5331 3398
rect -5293 3001 -5287 3398
rect -5337 2989 -5287 3001
rect -5171 3398 -5121 3410
rect -5171 3001 -5165 3398
rect -5127 3001 -5121 3398
rect -5171 2989 -5121 3001
rect -5005 3398 -4955 3410
rect -5005 3001 -4999 3398
rect -4961 3001 -4955 3398
rect -5005 2989 -4955 3001
rect -4839 3398 -4789 3410
rect -4839 3001 -4833 3398
rect -4795 3001 -4789 3398
rect -4839 2989 -4789 3001
rect -4673 3398 -4623 3410
rect -4673 3001 -4667 3398
rect -4629 3001 -4623 3398
rect -4673 2989 -4623 3001
rect -4507 3398 -4457 3410
rect -4507 3001 -4501 3398
rect -4463 3001 -4457 3398
rect -4507 2989 -4457 3001
rect -4341 3398 -4291 3410
rect -4341 3001 -4335 3398
rect -4297 3001 -4291 3398
rect -4341 2989 -4291 3001
rect -4175 3398 -4125 3410
rect -4175 3001 -4169 3398
rect -4131 3001 -4125 3398
rect -4175 2989 -4125 3001
rect -4009 3398 -3959 3410
rect -4009 3001 -4003 3398
rect -3965 3001 -3959 3398
rect -4009 2989 -3959 3001
rect -3843 3398 -3793 3410
rect -3843 3001 -3837 3398
rect -3799 3001 -3793 3398
rect -3843 2989 -3793 3001
rect -3677 3398 -3627 3410
rect -3677 3001 -3671 3398
rect -3633 3001 -3627 3398
rect -3677 2989 -3627 3001
rect -3511 3398 -3461 3410
rect -3511 3001 -3505 3398
rect -3467 3001 -3461 3398
rect -3511 2989 -3461 3001
rect -3345 3398 -3295 3410
rect -3345 3001 -3339 3398
rect -3301 3001 -3295 3398
rect -3345 2989 -3295 3001
rect -3179 3398 -3129 3410
rect -3179 3001 -3173 3398
rect -3135 3001 -3129 3398
rect -3179 2989 -3129 3001
rect -3013 3398 -2963 3410
rect -3013 3001 -3007 3398
rect -2969 3001 -2963 3398
rect -3013 2989 -2963 3001
rect -2847 3398 -2797 3410
rect -2847 3001 -2841 3398
rect -2803 3001 -2797 3398
rect -2847 2989 -2797 3001
rect -2681 3398 -2631 3410
rect -2681 3001 -2675 3398
rect -2637 3001 -2631 3398
rect -2681 2989 -2631 3001
rect -2515 3398 -2465 3410
rect -2515 3001 -2509 3398
rect -2471 3001 -2465 3398
rect -2515 2989 -2465 3001
rect -2349 3398 -2299 3410
rect -2349 3001 -2343 3398
rect -2305 3001 -2299 3398
rect -2349 2989 -2299 3001
rect -2183 3398 -2133 3410
rect -2183 3001 -2177 3398
rect -2139 3001 -2133 3398
rect -2183 2989 -2133 3001
rect -2017 3398 -1967 3410
rect -2017 3001 -2011 3398
rect -1973 3001 -1967 3398
rect -2017 2989 -1967 3001
rect -1851 3398 -1801 3410
rect -1851 3001 -1845 3398
rect -1807 3001 -1801 3398
rect -1851 2989 -1801 3001
rect -1685 3398 -1635 3410
rect -1685 3001 -1679 3398
rect -1641 3001 -1635 3398
rect -1685 2989 -1635 3001
rect -1519 3398 -1469 3410
rect -1519 3001 -1513 3398
rect -1475 3001 -1469 3398
rect -1519 2989 -1469 3001
rect -1353 3398 -1303 3410
rect -1353 3001 -1347 3398
rect -1309 3001 -1303 3398
rect -1353 2989 -1303 3001
rect -1187 3398 -1137 3410
rect -1187 3001 -1181 3398
rect -1143 3001 -1137 3398
rect -1187 2989 -1137 3001
rect -1021 3398 -971 3410
rect -1021 3001 -1015 3398
rect -977 3001 -971 3398
rect -1021 2989 -971 3001
rect -855 3398 -805 3410
rect -855 3001 -849 3398
rect -811 3001 -805 3398
rect -855 2989 -805 3001
rect -689 3398 -639 3410
rect -689 3001 -683 3398
rect -645 3001 -639 3398
rect -689 2989 -639 3001
rect -523 3398 -473 3410
rect -523 3001 -517 3398
rect -479 3001 -473 3398
rect -523 2989 -473 3001
rect -357 3398 -307 3410
rect -357 3001 -351 3398
rect -313 3001 -307 3398
rect -357 2989 -307 3001
rect -191 3398 -141 3410
rect -191 3001 -185 3398
rect -147 3001 -141 3398
rect -191 2989 -141 3001
rect -25 3398 25 3410
rect -25 3001 -19 3398
rect 19 3001 25 3398
rect -25 2989 25 3001
rect 141 3398 191 3410
rect 141 3001 147 3398
rect 185 3001 191 3398
rect 141 2989 191 3001
rect 307 3398 357 3410
rect 307 3001 313 3398
rect 351 3001 357 3398
rect 307 2989 357 3001
rect 473 3398 523 3410
rect 473 3001 479 3398
rect 517 3001 523 3398
rect 473 2989 523 3001
rect 639 3398 689 3410
rect 639 3001 645 3398
rect 683 3001 689 3398
rect 639 2989 689 3001
rect 805 3398 855 3410
rect 805 3001 811 3398
rect 849 3001 855 3398
rect 805 2989 855 3001
rect 971 3398 1021 3410
rect 971 3001 977 3398
rect 1015 3001 1021 3398
rect 971 2989 1021 3001
rect 1137 3398 1187 3410
rect 1137 3001 1143 3398
rect 1181 3001 1187 3398
rect 1137 2989 1187 3001
rect 1303 3398 1353 3410
rect 1303 3001 1309 3398
rect 1347 3001 1353 3398
rect 1303 2989 1353 3001
rect 1469 3398 1519 3410
rect 1469 3001 1475 3398
rect 1513 3001 1519 3398
rect 1469 2989 1519 3001
rect 1635 3398 1685 3410
rect 1635 3001 1641 3398
rect 1679 3001 1685 3398
rect 1635 2989 1685 3001
rect 1801 3398 1851 3410
rect 1801 3001 1807 3398
rect 1845 3001 1851 3398
rect 1801 2989 1851 3001
rect 1967 3398 2017 3410
rect 1967 3001 1973 3398
rect 2011 3001 2017 3398
rect 1967 2989 2017 3001
rect 2133 3398 2183 3410
rect 2133 3001 2139 3398
rect 2177 3001 2183 3398
rect 2133 2989 2183 3001
rect 2299 3398 2349 3410
rect 2299 3001 2305 3398
rect 2343 3001 2349 3398
rect 2299 2989 2349 3001
rect 2465 3398 2515 3410
rect 2465 3001 2471 3398
rect 2509 3001 2515 3398
rect 2465 2989 2515 3001
rect 2631 3398 2681 3410
rect 2631 3001 2637 3398
rect 2675 3001 2681 3398
rect 2631 2989 2681 3001
rect 2797 3398 2847 3410
rect 2797 3001 2803 3398
rect 2841 3001 2847 3398
rect 2797 2989 2847 3001
rect 2963 3398 3013 3410
rect 2963 3001 2969 3398
rect 3007 3001 3013 3398
rect 2963 2989 3013 3001
rect 3129 3398 3179 3410
rect 3129 3001 3135 3398
rect 3173 3001 3179 3398
rect 3129 2989 3179 3001
rect 3295 3398 3345 3410
rect 3295 3001 3301 3398
rect 3339 3001 3345 3398
rect 3295 2989 3345 3001
rect 3461 3398 3511 3410
rect 3461 3001 3467 3398
rect 3505 3001 3511 3398
rect 3461 2989 3511 3001
rect 3627 3398 3677 3410
rect 3627 3001 3633 3398
rect 3671 3001 3677 3398
rect 3627 2989 3677 3001
rect 3793 3398 3843 3410
rect 3793 3001 3799 3398
rect 3837 3001 3843 3398
rect 3793 2989 3843 3001
rect 3959 3398 4009 3410
rect 3959 3001 3965 3398
rect 4003 3001 4009 3398
rect 3959 2989 4009 3001
rect 4125 3398 4175 3410
rect 4125 3001 4131 3398
rect 4169 3001 4175 3398
rect 4125 2989 4175 3001
rect 4291 3398 4341 3410
rect 4291 3001 4297 3398
rect 4335 3001 4341 3398
rect 4291 2989 4341 3001
rect 4457 3398 4507 3410
rect 4457 3001 4463 3398
rect 4501 3001 4507 3398
rect 4457 2989 4507 3001
rect 4623 3398 4673 3410
rect 4623 3001 4629 3398
rect 4667 3001 4673 3398
rect 4623 2989 4673 3001
rect 4789 3398 4839 3410
rect 4789 3001 4795 3398
rect 4833 3001 4839 3398
rect 4789 2989 4839 3001
rect 4955 3398 5005 3410
rect 4955 3001 4961 3398
rect 4999 3001 5005 3398
rect 4955 2989 5005 3001
rect 5121 3398 5171 3410
rect 5121 3001 5127 3398
rect 5165 3001 5171 3398
rect 5121 2989 5171 3001
rect 5287 3398 5337 3410
rect 5287 3001 5293 3398
rect 5331 3001 5337 3398
rect 5287 2989 5337 3001
rect 5453 3398 5503 3410
rect 5453 3001 5459 3398
rect 5497 3001 5503 3398
rect 5453 2989 5503 3001
rect -5649 2810 -5603 2822
rect -5649 -2810 -5643 2810
rect -5609 -2810 -5603 2810
rect -5649 -2822 -5603 -2810
rect 5603 2810 5649 2822
rect 5603 -2810 5609 2810
rect 5643 -2810 5649 2810
rect 5603 -2822 5649 -2810
rect -5503 -3001 -5453 -2989
rect -5503 -3398 -5497 -3001
rect -5459 -3398 -5453 -3001
rect -5503 -3410 -5453 -3398
rect -5337 -3001 -5287 -2989
rect -5337 -3398 -5331 -3001
rect -5293 -3398 -5287 -3001
rect -5337 -3410 -5287 -3398
rect -5171 -3001 -5121 -2989
rect -5171 -3398 -5165 -3001
rect -5127 -3398 -5121 -3001
rect -5171 -3410 -5121 -3398
rect -5005 -3001 -4955 -2989
rect -5005 -3398 -4999 -3001
rect -4961 -3398 -4955 -3001
rect -5005 -3410 -4955 -3398
rect -4839 -3001 -4789 -2989
rect -4839 -3398 -4833 -3001
rect -4795 -3398 -4789 -3001
rect -4839 -3410 -4789 -3398
rect -4673 -3001 -4623 -2989
rect -4673 -3398 -4667 -3001
rect -4629 -3398 -4623 -3001
rect -4673 -3410 -4623 -3398
rect -4507 -3001 -4457 -2989
rect -4507 -3398 -4501 -3001
rect -4463 -3398 -4457 -3001
rect -4507 -3410 -4457 -3398
rect -4341 -3001 -4291 -2989
rect -4341 -3398 -4335 -3001
rect -4297 -3398 -4291 -3001
rect -4341 -3410 -4291 -3398
rect -4175 -3001 -4125 -2989
rect -4175 -3398 -4169 -3001
rect -4131 -3398 -4125 -3001
rect -4175 -3410 -4125 -3398
rect -4009 -3001 -3959 -2989
rect -4009 -3398 -4003 -3001
rect -3965 -3398 -3959 -3001
rect -4009 -3410 -3959 -3398
rect -3843 -3001 -3793 -2989
rect -3843 -3398 -3837 -3001
rect -3799 -3398 -3793 -3001
rect -3843 -3410 -3793 -3398
rect -3677 -3001 -3627 -2989
rect -3677 -3398 -3671 -3001
rect -3633 -3398 -3627 -3001
rect -3677 -3410 -3627 -3398
rect -3511 -3001 -3461 -2989
rect -3511 -3398 -3505 -3001
rect -3467 -3398 -3461 -3001
rect -3511 -3410 -3461 -3398
rect -3345 -3001 -3295 -2989
rect -3345 -3398 -3339 -3001
rect -3301 -3398 -3295 -3001
rect -3345 -3410 -3295 -3398
rect -3179 -3001 -3129 -2989
rect -3179 -3398 -3173 -3001
rect -3135 -3398 -3129 -3001
rect -3179 -3410 -3129 -3398
rect -3013 -3001 -2963 -2989
rect -3013 -3398 -3007 -3001
rect -2969 -3398 -2963 -3001
rect -3013 -3410 -2963 -3398
rect -2847 -3001 -2797 -2989
rect -2847 -3398 -2841 -3001
rect -2803 -3398 -2797 -3001
rect -2847 -3410 -2797 -3398
rect -2681 -3001 -2631 -2989
rect -2681 -3398 -2675 -3001
rect -2637 -3398 -2631 -3001
rect -2681 -3410 -2631 -3398
rect -2515 -3001 -2465 -2989
rect -2515 -3398 -2509 -3001
rect -2471 -3398 -2465 -3001
rect -2515 -3410 -2465 -3398
rect -2349 -3001 -2299 -2989
rect -2349 -3398 -2343 -3001
rect -2305 -3398 -2299 -3001
rect -2349 -3410 -2299 -3398
rect -2183 -3001 -2133 -2989
rect -2183 -3398 -2177 -3001
rect -2139 -3398 -2133 -3001
rect -2183 -3410 -2133 -3398
rect -2017 -3001 -1967 -2989
rect -2017 -3398 -2011 -3001
rect -1973 -3398 -1967 -3001
rect -2017 -3410 -1967 -3398
rect -1851 -3001 -1801 -2989
rect -1851 -3398 -1845 -3001
rect -1807 -3398 -1801 -3001
rect -1851 -3410 -1801 -3398
rect -1685 -3001 -1635 -2989
rect -1685 -3398 -1679 -3001
rect -1641 -3398 -1635 -3001
rect -1685 -3410 -1635 -3398
rect -1519 -3001 -1469 -2989
rect -1519 -3398 -1513 -3001
rect -1475 -3398 -1469 -3001
rect -1519 -3410 -1469 -3398
rect -1353 -3001 -1303 -2989
rect -1353 -3398 -1347 -3001
rect -1309 -3398 -1303 -3001
rect -1353 -3410 -1303 -3398
rect -1187 -3001 -1137 -2989
rect -1187 -3398 -1181 -3001
rect -1143 -3398 -1137 -3001
rect -1187 -3410 -1137 -3398
rect -1021 -3001 -971 -2989
rect -1021 -3398 -1015 -3001
rect -977 -3398 -971 -3001
rect -1021 -3410 -971 -3398
rect -855 -3001 -805 -2989
rect -855 -3398 -849 -3001
rect -811 -3398 -805 -3001
rect -855 -3410 -805 -3398
rect -689 -3001 -639 -2989
rect -689 -3398 -683 -3001
rect -645 -3398 -639 -3001
rect -689 -3410 -639 -3398
rect -523 -3001 -473 -2989
rect -523 -3398 -517 -3001
rect -479 -3398 -473 -3001
rect -523 -3410 -473 -3398
rect -357 -3001 -307 -2989
rect -357 -3398 -351 -3001
rect -313 -3398 -307 -3001
rect -357 -3410 -307 -3398
rect -191 -3001 -141 -2989
rect -191 -3398 -185 -3001
rect -147 -3398 -141 -3001
rect -191 -3410 -141 -3398
rect -25 -3001 25 -2989
rect -25 -3398 -19 -3001
rect 19 -3398 25 -3001
rect -25 -3410 25 -3398
rect 141 -3001 191 -2989
rect 141 -3398 147 -3001
rect 185 -3398 191 -3001
rect 141 -3410 191 -3398
rect 307 -3001 357 -2989
rect 307 -3398 313 -3001
rect 351 -3398 357 -3001
rect 307 -3410 357 -3398
rect 473 -3001 523 -2989
rect 473 -3398 479 -3001
rect 517 -3398 523 -3001
rect 473 -3410 523 -3398
rect 639 -3001 689 -2989
rect 639 -3398 645 -3001
rect 683 -3398 689 -3001
rect 639 -3410 689 -3398
rect 805 -3001 855 -2989
rect 805 -3398 811 -3001
rect 849 -3398 855 -3001
rect 805 -3410 855 -3398
rect 971 -3001 1021 -2989
rect 971 -3398 977 -3001
rect 1015 -3398 1021 -3001
rect 971 -3410 1021 -3398
rect 1137 -3001 1187 -2989
rect 1137 -3398 1143 -3001
rect 1181 -3398 1187 -3001
rect 1137 -3410 1187 -3398
rect 1303 -3001 1353 -2989
rect 1303 -3398 1309 -3001
rect 1347 -3398 1353 -3001
rect 1303 -3410 1353 -3398
rect 1469 -3001 1519 -2989
rect 1469 -3398 1475 -3001
rect 1513 -3398 1519 -3001
rect 1469 -3410 1519 -3398
rect 1635 -3001 1685 -2989
rect 1635 -3398 1641 -3001
rect 1679 -3398 1685 -3001
rect 1635 -3410 1685 -3398
rect 1801 -3001 1851 -2989
rect 1801 -3398 1807 -3001
rect 1845 -3398 1851 -3001
rect 1801 -3410 1851 -3398
rect 1967 -3001 2017 -2989
rect 1967 -3398 1973 -3001
rect 2011 -3398 2017 -3001
rect 1967 -3410 2017 -3398
rect 2133 -3001 2183 -2989
rect 2133 -3398 2139 -3001
rect 2177 -3398 2183 -3001
rect 2133 -3410 2183 -3398
rect 2299 -3001 2349 -2989
rect 2299 -3398 2305 -3001
rect 2343 -3398 2349 -3001
rect 2299 -3410 2349 -3398
rect 2465 -3001 2515 -2989
rect 2465 -3398 2471 -3001
rect 2509 -3398 2515 -3001
rect 2465 -3410 2515 -3398
rect 2631 -3001 2681 -2989
rect 2631 -3398 2637 -3001
rect 2675 -3398 2681 -3001
rect 2631 -3410 2681 -3398
rect 2797 -3001 2847 -2989
rect 2797 -3398 2803 -3001
rect 2841 -3398 2847 -3001
rect 2797 -3410 2847 -3398
rect 2963 -3001 3013 -2989
rect 2963 -3398 2969 -3001
rect 3007 -3398 3013 -3001
rect 2963 -3410 3013 -3398
rect 3129 -3001 3179 -2989
rect 3129 -3398 3135 -3001
rect 3173 -3398 3179 -3001
rect 3129 -3410 3179 -3398
rect 3295 -3001 3345 -2989
rect 3295 -3398 3301 -3001
rect 3339 -3398 3345 -3001
rect 3295 -3410 3345 -3398
rect 3461 -3001 3511 -2989
rect 3461 -3398 3467 -3001
rect 3505 -3398 3511 -3001
rect 3461 -3410 3511 -3398
rect 3627 -3001 3677 -2989
rect 3627 -3398 3633 -3001
rect 3671 -3398 3677 -3001
rect 3627 -3410 3677 -3398
rect 3793 -3001 3843 -2989
rect 3793 -3398 3799 -3001
rect 3837 -3398 3843 -3001
rect 3793 -3410 3843 -3398
rect 3959 -3001 4009 -2989
rect 3959 -3398 3965 -3001
rect 4003 -3398 4009 -3001
rect 3959 -3410 4009 -3398
rect 4125 -3001 4175 -2989
rect 4125 -3398 4131 -3001
rect 4169 -3398 4175 -3001
rect 4125 -3410 4175 -3398
rect 4291 -3001 4341 -2989
rect 4291 -3398 4297 -3001
rect 4335 -3398 4341 -3001
rect 4291 -3410 4341 -3398
rect 4457 -3001 4507 -2989
rect 4457 -3398 4463 -3001
rect 4501 -3398 4507 -3001
rect 4457 -3410 4507 -3398
rect 4623 -3001 4673 -2989
rect 4623 -3398 4629 -3001
rect 4667 -3398 4673 -3001
rect 4623 -3410 4673 -3398
rect 4789 -3001 4839 -2989
rect 4789 -3398 4795 -3001
rect 4833 -3398 4839 -3001
rect 4789 -3410 4839 -3398
rect 4955 -3001 5005 -2989
rect 4955 -3398 4961 -3001
rect 4999 -3398 5005 -3001
rect 4955 -3410 5005 -3398
rect 5121 -3001 5171 -2989
rect 5121 -3398 5127 -3001
rect 5165 -3398 5171 -3001
rect 5121 -3410 5171 -3398
rect 5287 -3001 5337 -2989
rect 5287 -3398 5293 -3001
rect 5331 -3398 5337 -3001
rect 5287 -3410 5337 -3398
rect 5453 -3001 5503 -2989
rect 5453 -3398 5459 -3001
rect 5497 -3398 5503 -3001
rect 5453 -3410 5503 -3398
rect -5621 -3512 5621 -3506
rect -5621 -3546 -5609 -3512
rect 5609 -3546 5621 -3512
rect -5621 -3552 5621 -3546
<< properties >>
string FIXED_BBOX -5626 -3529 5626 3529
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 30 m 1 nx 67 wmin 0.350 lmin 0.50 rho 319.8 val 28.524k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 100 viagt 100 viagl 80 viagr 80
<< end >>
