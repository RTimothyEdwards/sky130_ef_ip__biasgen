magic
tech sky130A
magscale 1 2
timestamp 1747752771
<< error_s >>
rect 134998 -2835 135078 -2549
rect 134998 -9375 135284 -2835
rect 134998 -10275 135978 -9375
rect 134998 -10561 135078 -10275
<< dnwell >>
rect 96152 17373 138230 25225
rect 89743 7999 138229 15851
rect 89743 -1114 138229 6738
rect 135078 -10481 138229 -2629
<< nwell >>
rect 96043 25019 138339 25334
rect 96043 17579 96358 25019
rect 138024 17579 138339 25019
rect 96043 17264 138339 17579
rect 89634 15645 138338 15960
rect 89634 8205 89949 15645
rect 138023 8205 138338 15645
rect 89634 7890 138338 8205
rect 89634 6532 138338 6847
rect 89634 -908 89949 6532
rect 138023 -908 138338 6532
rect 89634 -1223 138338 -908
rect 135078 -2835 138338 -2520
rect 138023 -10275 138338 -2835
rect 135078 -10590 138338 -10275
<< pwell >>
rect 125398 24997 125486 25019
rect 108895 8205 108983 8227
rect 108895 6510 108983 6532
<< mvpsubdiff >>
rect 95923 25446 95983 25480
rect 137413 25446 137603 25480
rect 138399 25446 138459 25480
rect 95923 25420 95957 25446
rect 88537 24692 88597 24726
rect 95249 24692 95309 24726
rect 88537 24666 95309 24692
rect 88571 24598 95275 24666
rect 88571 24503 88680 24598
rect 95204 24503 95275 24598
rect 88571 24469 89596 24503
rect 94944 24469 95275 24503
rect 88571 22875 88680 24469
rect 95204 22875 95275 24469
rect 88571 22841 89596 22875
rect 94944 22841 95275 22875
rect 88571 21247 88680 22841
rect 95204 21247 95275 22841
rect 88571 21213 89596 21247
rect 94944 21213 95275 21247
rect 88571 19619 88680 21213
rect 95204 19619 95275 21213
rect 88571 19585 89596 19619
rect 94944 19585 95275 19619
rect 88571 17991 88680 19585
rect 95204 17991 95275 19585
rect 88571 17957 89596 17991
rect 94944 17957 95275 17991
rect 88571 17856 88680 17957
rect 95204 17856 95275 17957
rect 88571 17788 95275 17856
rect 88537 17762 95309 17788
rect 88537 17728 88597 17762
rect 95249 17728 95309 17762
rect 138425 25420 138459 25446
rect 95923 17174 95957 17200
rect 138425 17174 138459 17200
rect 95923 17140 95983 17174
rect 137413 17140 137603 17174
rect 138399 17140 138459 17174
rect 89514 16050 89574 16084
rect 90370 16050 90560 16084
rect 138398 16050 138458 16084
rect 89514 16024 89548 16050
rect 138424 16024 138458 16050
rect 89514 7778 89548 7804
rect 138424 7778 138458 7804
rect 89514 7744 89574 7778
rect 138398 7744 138458 7778
rect 89514 6959 89574 6993
rect 90370 6959 90560 6993
rect 138398 6959 138458 6993
rect 89514 6933 89548 6959
rect 138424 6933 138458 6959
rect 89514 -1313 89548 -1287
rect 138424 -1313 138458 -1287
rect 89514 -1347 89574 -1313
rect 90370 -1347 90560 -1313
rect 138398 -1347 138458 -1313
rect 135144 -2430 135416 -2396
rect 138398 -2430 138458 -2396
rect 138424 -2456 138458 -2430
rect 138424 -10702 138458 -10676
rect 135144 -10736 135416 -10702
rect 138398 -10736 138458 -10702
<< mvnsubdiff >>
rect 96109 25248 138273 25268
rect 96109 25214 96189 25248
rect 137413 25214 137603 25248
rect 138193 25214 138273 25248
rect 96109 25194 138273 25214
rect 96109 25188 96183 25194
rect 96109 17410 96129 25188
rect 96163 17410 96183 25188
rect 96109 17404 96183 17410
rect 138199 25188 138273 25194
rect 138199 17410 138219 25188
rect 138253 17410 138273 25188
rect 138199 17404 138273 17410
rect 96109 17384 138273 17404
rect 96109 17350 96189 17384
rect 137413 17350 137603 17384
rect 138193 17350 138273 17384
rect 96109 17330 138273 17350
rect 89700 15874 138272 15894
rect 89700 15840 89780 15874
rect 90370 15840 90560 15874
rect 138192 15840 138272 15874
rect 89700 15820 138272 15840
rect 89700 15814 89774 15820
rect 89700 8036 89720 15814
rect 89754 8036 89774 15814
rect 89700 8030 89774 8036
rect 138198 15814 138272 15820
rect 138198 8036 138218 15814
rect 138252 8036 138272 15814
rect 138198 8030 138272 8036
rect 89700 8010 138272 8030
rect 89700 7976 89780 8010
rect 90370 7976 90560 8010
rect 138192 7976 138272 8010
rect 89700 7956 138272 7976
rect 89700 6761 138272 6781
rect 89700 6727 89780 6761
rect 90370 6727 90560 6761
rect 138192 6727 138272 6761
rect 89700 6707 138272 6727
rect 89700 6701 89774 6707
rect 89700 -1077 89720 6701
rect 89754 -1077 89774 6701
rect 89700 -1083 89774 -1077
rect 138198 6701 138272 6707
rect 138198 -1077 138218 6701
rect 138252 -1077 138272 6701
rect 138198 -1083 138272 -1077
rect 89700 -1103 138272 -1083
rect 89700 -1137 89780 -1103
rect 90370 -1137 90560 -1103
rect 138192 -1137 138272 -1103
rect 89700 -1157 138272 -1137
rect 135144 -2606 138272 -2586
rect 135144 -2640 135416 -2606
rect 138192 -2640 138272 -2606
rect 135144 -2660 138272 -2640
rect 138198 -2666 138272 -2660
rect 138198 -10444 138218 -2666
rect 138252 -10444 138272 -2666
rect 138198 -10450 138272 -10444
rect 135144 -10470 138272 -10450
rect 135144 -10504 135416 -10470
rect 138192 -10504 138272 -10470
rect 135144 -10524 138272 -10504
<< mvpsubdiffcont >>
rect 95983 25446 137413 25480
rect 137603 25446 138399 25480
rect 88597 24692 95249 24726
rect 88537 17788 88571 24666
rect 95275 17788 95309 24666
rect 88597 17728 95249 17762
rect 95923 17200 95957 25420
rect 138425 17200 138459 25420
rect 95983 17140 137413 17174
rect 137603 17140 138399 17174
rect 89574 16050 90370 16084
rect 90560 16050 138398 16084
rect 89514 7804 89548 16024
rect 138424 7804 138458 16024
rect 89574 7744 138398 7778
rect 89574 6959 90370 6993
rect 90560 6959 138398 6993
rect 89514 -1287 89548 6933
rect 138424 -1287 138458 6933
rect 89574 -1347 90370 -1313
rect 90560 -1347 138398 -1313
rect 135416 -2430 138398 -2396
rect 138424 -10676 138458 -2456
rect 135416 -10736 138398 -10702
<< mvnsubdiffcont >>
rect 96189 25214 137413 25248
rect 137603 25214 138193 25248
rect 96129 17410 96163 25188
rect 138219 17410 138253 25188
rect 96189 17350 137413 17384
rect 137603 17350 138193 17384
rect 89780 15840 90370 15874
rect 90560 15840 138192 15874
rect 89720 8036 89754 15814
rect 138218 8036 138252 15814
rect 89780 7976 90370 8010
rect 90560 7976 138192 8010
rect 89780 6727 90370 6761
rect 90560 6727 138192 6761
rect 89720 -1077 89754 6701
rect 138218 -1077 138252 6701
rect 89780 -1137 90370 -1103
rect 90560 -1137 138192 -1103
rect 135416 -2640 138192 -2606
rect 138218 -10444 138252 -2666
rect 135416 -10504 138192 -10470
<< locali >>
rect 95923 25446 95983 25480
rect 95923 25430 96074 25446
rect 95923 25420 95969 25430
rect 95220 24726 95923 24727
rect 88537 24692 88597 24726
rect 95249 24692 95923 24726
rect 88537 24666 95923 24692
rect 88571 24604 95275 24666
rect 88571 17850 88665 24604
rect 90110 24164 90280 24180
rect 90110 24062 90131 24164
rect 90264 24062 90280 24164
rect 90110 24046 90280 24062
rect 92702 24164 92872 24180
rect 92702 24062 92723 24164
rect 92856 24062 92872 24164
rect 92702 24046 92872 24062
rect 91871 23168 91918 23234
rect 94456 23170 94557 23235
rect 90110 22536 90280 22552
rect 90110 22434 90131 22536
rect 90264 22434 90280 22536
rect 90110 22418 90280 22434
rect 92702 22536 92872 22552
rect 92702 22434 92723 22536
rect 92856 22434 92872 22536
rect 92702 22418 92872 22434
rect 91871 21540 91918 21606
rect 94444 21542 94545 21607
rect 90110 20908 90280 20924
rect 90110 20806 90131 20908
rect 90264 20806 90280 20908
rect 90110 20790 90280 20806
rect 92702 20908 92872 20924
rect 92702 20806 92723 20908
rect 92856 20806 92872 20908
rect 92702 20790 92872 20806
rect 91871 20047 91879 20087
rect 91871 19912 91918 19978
rect 94453 19910 94554 19975
rect 90110 19280 90280 19296
rect 90110 19178 90131 19280
rect 90264 19178 90280 19280
rect 90110 19162 90280 19178
rect 92702 19280 92872 19296
rect 92702 19178 92723 19280
rect 92856 19178 92872 19280
rect 92702 19162 92872 19178
rect 91871 18416 91879 18456
rect 91871 18284 91918 18350
rect 94444 18285 94545 18350
rect 95192 17850 95275 24604
rect 88571 17788 95275 17850
rect 95309 24530 95923 24666
rect 95309 17788 95923 17925
rect 88537 17762 95923 17788
rect 88537 17728 88597 17762
rect 95249 17728 95923 17762
rect 95957 17200 95969 25420
rect 95923 17189 95969 17200
rect 96021 25421 96074 25430
rect 137413 25421 137603 25480
rect 138399 25446 138459 25480
rect 138308 25430 138459 25446
rect 138308 25421 138361 25430
rect 96021 25334 138361 25421
rect 96021 17273 96065 25334
rect 96129 25214 96189 25248
rect 137413 25214 137603 25248
rect 138193 25214 138253 25248
rect 96129 25192 138253 25214
rect 96129 25188 96194 25192
rect 96163 17415 96194 25188
rect 96253 25035 138129 25192
rect 96253 17569 96300 25035
rect 138082 17569 138129 25035
rect 96253 17415 138129 17569
rect 138188 25188 138253 25192
rect 138188 17415 138219 25188
rect 96163 17410 138219 17415
rect 96129 17384 138253 17410
rect 96129 17350 96189 17384
rect 137413 17350 137603 17384
rect 138193 17350 138253 17384
rect 138317 17273 138361 25334
rect 96021 17189 138361 17273
rect 138413 25420 138459 25430
rect 138413 17200 138425 25420
rect 138459 24530 138541 24727
rect 138413 17189 138459 17200
rect 95923 17174 138459 17189
rect 95923 17140 95983 17174
rect 137413 17140 137603 17174
rect 138399 17140 138459 17174
rect 89514 16050 89574 16084
rect 90370 16050 90560 16084
rect 138398 16050 138458 16084
rect 89514 16035 138458 16050
rect 89514 16024 89560 16035
rect 89432 8497 89514 8694
rect 89548 7804 89560 16024
rect 89514 7794 89560 7804
rect 89612 15951 138360 16035
rect 89612 7890 89656 15951
rect 89720 15840 89780 15874
rect 90370 15840 90560 15874
rect 138192 15840 138252 15874
rect 89720 15814 138252 15840
rect 89754 15809 138218 15814
rect 89754 8036 89785 15809
rect 89720 8032 89785 8036
rect 89844 15655 138128 15809
rect 89844 8189 89891 15655
rect 90874 15549 90993 15655
rect 138081 8189 138128 15655
rect 89844 8032 138128 8189
rect 138187 8036 138218 15809
rect 138187 8032 138252 8036
rect 89720 8010 138252 8032
rect 89720 7976 89780 8010
rect 90370 7976 90560 8010
rect 138192 7976 138252 8010
rect 138316 7890 138360 15951
rect 89612 7803 138360 7890
rect 89612 7794 89665 7803
rect 89514 7778 89665 7794
rect 138307 7794 138360 7803
rect 138412 16024 138458 16035
rect 138412 7804 138424 16024
rect 138458 8497 138540 8694
rect 138412 7794 138458 7804
rect 138307 7778 138458 7794
rect 89514 7744 89574 7778
rect 138398 7744 138458 7778
rect 89514 6959 89574 6993
rect 89514 6943 89665 6959
rect 89514 6933 89560 6943
rect 89432 6043 89514 6240
rect 89548 -1287 89560 6933
rect 89514 -1298 89560 -1287
rect 89612 6934 89665 6943
rect 90370 6934 90560 6993
rect 138398 6959 138458 6993
rect 138307 6943 138458 6959
rect 138307 6934 138360 6943
rect 89612 6847 138360 6934
rect 89612 -1214 89656 6847
rect 89720 6727 89780 6761
rect 90370 6727 90560 6761
rect 138192 6727 138252 6761
rect 89720 6705 138252 6727
rect 89720 6701 89785 6705
rect 89754 -1072 89785 6701
rect 89844 6548 138128 6705
rect 89844 -918 89891 6548
rect 138081 -918 138128 6548
rect 89844 -1072 138128 -918
rect 138187 6701 138252 6705
rect 138187 -1072 138218 6701
rect 89754 -1077 138218 -1072
rect 89720 -1103 138252 -1077
rect 89720 -1137 89780 -1103
rect 90370 -1137 90560 -1103
rect 138192 -1137 138252 -1103
rect 138316 -1214 138360 6847
rect 89612 -1298 138360 -1214
rect 138412 6933 138458 6943
rect 138412 -1287 138424 6933
rect 138458 6043 138540 6240
rect 138412 -1298 138458 -1287
rect 89514 -1313 138458 -1298
rect 89514 -1347 89574 -1313
rect 90370 -1347 90560 -1313
rect 138398 -1347 138458 -1313
rect 135144 -2430 135416 -2396
rect 138398 -2430 138458 -2396
rect 135144 -2445 138458 -2430
rect 135144 -2529 138360 -2445
rect 135152 -2640 135416 -2606
rect 138192 -2640 138252 -2606
rect 135152 -2666 138252 -2640
rect 135152 -2671 138218 -2666
rect 135152 -2825 138128 -2671
rect 138081 -10291 138128 -2825
rect 135144 -10448 138128 -10291
rect 138187 -10444 138218 -2671
rect 138187 -10448 138252 -10444
rect 135144 -10470 138252 -10448
rect 135144 -10504 135416 -10470
rect 138192 -10504 138252 -10470
rect 138316 -10590 138360 -2529
rect 135144 -10677 138360 -10590
rect 135144 -10736 135416 -10677
rect 138307 -10686 138360 -10677
rect 138412 -2456 138458 -2445
rect 138412 -10676 138424 -2456
rect 138458 -9983 138540 -9786
rect 138412 -10686 138458 -10676
rect 138307 -10702 138458 -10686
rect 138398 -10736 138458 -10702
<< viali >>
rect 96074 25446 137413 25465
rect 89666 24024 89702 24153
rect 90131 24062 90264 24164
rect 92723 24062 92856 24164
rect 89666 23224 89702 23353
rect 91823 23281 91871 23512
rect 94415 23281 94463 23512
rect 92206 23025 92252 23204
rect 94798 23025 94844 23204
rect 89666 22396 89702 22525
rect 90131 22434 90264 22536
rect 92723 22434 92856 22536
rect 89666 21596 89702 21725
rect 91823 21653 91871 21884
rect 94415 21653 94463 21884
rect 92206 21397 92252 21576
rect 94798 21397 94844 21576
rect 89666 20768 89702 20897
rect 90131 20806 90264 20908
rect 92723 20806 92856 20908
rect 89666 19968 89702 20097
rect 91823 20025 91871 20256
rect 94415 20025 94463 20256
rect 92206 19769 92252 19948
rect 94798 19769 94844 19948
rect 89666 19140 89702 19269
rect 90131 19178 90264 19280
rect 92723 19178 92856 19280
rect 89666 18340 89702 18469
rect 91823 18397 91871 18628
rect 94415 18397 94463 18628
rect 92206 18141 92252 18320
rect 94798 18141 94844 18320
rect 95969 17189 96021 25430
rect 96074 25421 137413 25446
rect 137603 25446 138308 25465
rect 137603 25421 138308 25446
rect 96194 17415 96253 25192
rect 138129 17415 138188 25192
rect 138361 17189 138413 25430
rect 89560 7794 89612 16035
rect 89785 8032 89844 15809
rect 90874 15439 90993 15549
rect 138128 8032 138187 15809
rect 89665 7778 138307 7803
rect 138360 7794 138412 16035
rect 89665 7759 138307 7778
rect 89665 6959 90370 6978
rect 89560 -1298 89612 6943
rect 89665 6934 90370 6959
rect 90560 6959 138307 6978
rect 90560 6934 138307 6959
rect 89785 -1072 89844 6705
rect 138128 -1072 138187 6705
rect 138360 -1298 138412 6943
rect 138128 -10448 138187 -2671
rect 135416 -10702 138307 -10677
rect 138360 -10686 138412 -2445
rect 135416 -10721 138307 -10702
<< metal1 >>
rect 95933 25465 138449 25480
rect 95933 25430 96074 25465
rect 95933 24634 95969 25430
rect 95759 24602 95969 24634
rect 96021 25421 96074 25430
rect 137413 25421 137603 25465
rect 138308 25430 138449 25465
rect 138308 25421 138361 25430
rect 96021 25402 138361 25421
rect 88825 24405 93088 24483
rect 94360 24405 95047 24483
rect 89654 24153 89714 24165
rect 89654 24024 89666 24153
rect 89702 24138 89714 24153
rect 90110 24164 90280 24180
rect 90110 24138 90131 24164
rect 89702 24088 90131 24138
rect 89702 24024 89714 24088
rect 90110 24062 90131 24088
rect 90264 24062 90280 24164
rect 90110 24046 90280 24062
rect 92702 24164 92872 24180
rect 92702 24062 92723 24164
rect 92856 24062 92872 24164
rect 92702 24046 92872 24062
rect 89654 24012 89714 24024
rect 89111 23825 89122 23882
rect 89505 23825 95047 23882
rect 88747 23588 90501 23761
rect 91780 23588 95047 23761
rect 91787 23547 91890 23551
rect 91810 23512 91883 23518
rect 89654 23353 89714 23365
rect 89654 23224 89666 23353
rect 89702 23224 89714 23353
rect 91810 23281 91823 23512
rect 91871 23498 91883 23512
rect 94402 23512 94475 23518
rect 91871 23494 91941 23498
rect 91871 23443 93852 23494
rect 91871 23298 91941 23443
rect 92690 23328 92696 23334
rect 91871 23281 91883 23298
rect 91810 23275 91883 23281
rect 92030 23288 92696 23328
rect 91826 23268 91866 23275
rect 89654 23220 89714 23224
rect 92030 23220 92070 23288
rect 92690 23282 92696 23288
rect 92748 23282 92754 23334
rect 89654 23212 92070 23220
rect 92200 23214 92259 23216
rect 89656 23180 92070 23212
rect 92199 23204 92207 23214
rect 92199 23025 92206 23204
rect 92259 23084 92265 23214
rect 93801 23183 93852 23443
rect 94402 23281 94415 23512
rect 94463 23444 94475 23512
rect 95385 23444 95391 23604
rect 94463 23404 95391 23444
rect 95443 23404 95449 23604
rect 95759 23463 95788 24602
rect 95759 23432 95969 23463
rect 94463 23281 94475 23404
rect 95734 23321 95740 23327
rect 94402 23275 94475 23281
rect 94418 23268 94458 23275
rect 94565 23270 95740 23321
rect 94565 23183 94616 23270
rect 93801 23132 94616 23183
rect 94789 23214 94852 23230
rect 92199 23014 92207 23025
rect 92259 23014 92265 23044
rect 94789 23014 94795 23214
rect 94847 23186 94852 23214
rect 94847 23014 94853 23186
rect 95734 23127 95740 23270
rect 95792 23127 95798 23327
rect 92199 23012 92265 23014
rect 94792 23013 94851 23014
rect 88791 22771 93083 22944
rect 94353 22771 95047 22944
rect 89654 22525 89714 22537
rect 89654 22396 89666 22525
rect 89702 22508 89714 22525
rect 90110 22536 90280 22552
rect 90110 22508 90131 22536
rect 89702 22458 90131 22508
rect 89702 22396 89714 22458
rect 90110 22434 90131 22458
rect 90264 22434 90280 22536
rect 90110 22418 90280 22434
rect 92702 22536 92872 22552
rect 92702 22434 92723 22536
rect 92856 22434 92872 22536
rect 92702 22418 92872 22434
rect 89654 22384 89714 22396
rect 89111 22197 89122 22254
rect 89505 22197 95047 22254
rect 88758 21949 90501 22122
rect 91780 21949 95047 22122
rect 91807 21886 91883 21890
rect 91807 21884 91939 21886
rect 89654 21725 89714 21737
rect 89654 21596 89666 21725
rect 89702 21596 89714 21725
rect 91807 21653 91823 21884
rect 91871 21883 91939 21884
rect 94399 21884 94475 21890
rect 91871 21832 94098 21883
rect 91871 21686 91939 21832
rect 92734 21717 92740 21723
rect 91871 21653 91883 21686
rect 91807 21647 91883 21653
rect 92014 21677 92740 21717
rect 91822 21643 91862 21647
rect 89654 21585 89714 21596
rect 92014 21585 92054 21677
rect 92734 21671 92740 21677
rect 92792 21671 92798 21723
rect 89654 21584 92054 21585
rect 89656 21545 92054 21584
rect 92200 21586 92259 21588
rect 92200 21576 92207 21586
rect 92200 21397 92206 21576
rect 92259 21456 92265 21586
rect 94047 21580 94098 21832
rect 94399 21653 94415 21884
rect 94463 21816 94475 21884
rect 95475 21816 95481 21976
rect 94463 21776 95481 21816
rect 95533 21816 95539 21976
rect 95713 21816 95719 21976
rect 95533 21776 95719 21816
rect 95771 21776 95777 21976
rect 94463 21653 94475 21776
rect 95556 21708 95651 21715
rect 94399 21647 94475 21653
rect 94584 21700 95651 21708
rect 94584 21693 95593 21700
rect 94584 21657 95060 21693
rect 94414 21643 94454 21647
rect 94584 21580 94635 21657
rect 94047 21529 94635 21580
rect 94782 21586 94852 21616
rect 94782 21576 94795 21586
rect 92200 21386 92207 21397
rect 92259 21386 92265 21416
rect 94789 21386 94795 21576
rect 94847 21555 94852 21586
rect 94847 21386 94853 21555
rect 95054 21493 95060 21657
rect 95112 21657 95593 21693
rect 95112 21493 95118 21657
rect 95587 21500 95593 21657
rect 95645 21500 95651 21700
rect 92200 21385 92265 21386
rect 94792 21385 94851 21386
rect 92201 21384 92265 21385
rect 88775 21149 93087 21322
rect 94357 21149 95047 21322
rect 89654 20897 89714 20909
rect 89654 20768 89666 20897
rect 89702 20880 89714 20897
rect 90110 20908 90280 20924
rect 90110 20880 90131 20908
rect 89702 20830 90131 20880
rect 89702 20768 89714 20830
rect 90110 20806 90131 20830
rect 90264 20806 90280 20908
rect 90110 20790 90280 20806
rect 92702 20908 92872 20924
rect 92702 20806 92723 20908
rect 92856 20806 92872 20908
rect 92702 20790 92872 20806
rect 89654 20756 89714 20768
rect 89111 20569 89125 20626
rect 89505 20569 95047 20626
rect 88747 20333 90505 20506
rect 91784 20333 95047 20506
rect 91807 20256 91883 20262
rect 89654 20097 89714 20109
rect 89654 19968 89666 20097
rect 89702 19970 89714 20097
rect 91807 20025 91823 20256
rect 91871 20247 91883 20256
rect 94399 20256 94475 20262
rect 91871 20244 91947 20247
rect 91871 20193 94149 20244
rect 91871 20047 91947 20193
rect 92724 20130 92730 20136
rect 92043 20090 92730 20130
rect 91871 20025 91883 20047
rect 91807 20019 91883 20025
rect 91822 20014 91862 20019
rect 92043 19970 92083 20090
rect 92724 20084 92730 20090
rect 92782 20084 92788 20136
rect 89702 19968 92083 19970
rect 89654 19930 92083 19968
rect 92201 19960 92241 19967
rect 94098 19962 94149 20193
rect 94399 20025 94415 20256
rect 94463 20188 94475 20256
rect 95557 20188 95563 20348
rect 94463 20148 95563 20188
rect 95615 20148 95621 20348
rect 94463 20025 94475 20148
rect 94399 20019 94475 20025
rect 94535 20056 95214 20072
rect 94535 20021 95183 20056
rect 94414 20014 94454 20019
rect 94535 19962 94586 20021
rect 92200 19958 92259 19960
rect 92199 19948 92207 19958
rect 92199 19769 92206 19948
rect 92199 19758 92207 19769
rect 92259 19758 92265 19958
rect 94098 19911 94586 19962
rect 94782 19958 94855 19988
rect 94782 19948 94795 19958
rect 94847 19948 94855 19958
rect 94789 19758 94795 19948
rect 94847 19758 94853 19948
rect 95177 19896 95183 20021
rect 95171 19856 95183 19896
rect 95235 19856 95241 20056
rect 92199 19756 92265 19758
rect 94792 19757 94851 19758
rect 88764 19522 93085 19695
rect 94355 19522 95047 19695
rect 89654 19269 89714 19281
rect 89654 19140 89666 19269
rect 89702 19248 89714 19269
rect 90110 19280 90280 19296
rect 90110 19248 90131 19280
rect 89702 19198 90131 19248
rect 89702 19140 89714 19198
rect 90110 19178 90131 19198
rect 90264 19178 90280 19280
rect 90110 19162 90280 19178
rect 92702 19280 92872 19296
rect 92702 19178 92723 19280
rect 92856 19178 92872 19280
rect 92702 19162 92872 19178
rect 89654 19128 89714 19140
rect 89111 18941 89129 18998
rect 89505 18941 95047 18998
rect 88764 18705 90501 18878
rect 91780 18705 95047 18878
rect 91807 18628 91883 18634
rect 89654 18469 89714 18481
rect 89654 18340 89666 18469
rect 89702 18340 89714 18469
rect 91807 18397 91823 18628
rect 91871 18616 91883 18628
rect 94399 18628 94475 18634
rect 91871 18613 91947 18616
rect 91871 18562 93749 18613
rect 91871 18416 91947 18562
rect 92693 18479 92699 18485
rect 92004 18439 92699 18479
rect 91871 18397 91883 18416
rect 91807 18391 91883 18397
rect 91822 18384 91862 18391
rect 89654 18335 89714 18340
rect 92004 18335 92044 18439
rect 92693 18433 92699 18439
rect 92751 18433 92757 18485
rect 89654 18328 92044 18335
rect 92201 18332 92241 18341
rect 89656 18295 92044 18328
rect 92200 18330 92259 18332
rect 92200 18320 92207 18330
rect 92200 18141 92206 18320
rect 92200 18130 92207 18141
rect 92259 18130 92265 18330
rect 93698 18279 93749 18562
rect 94399 18397 94415 18628
rect 94463 18560 94475 18628
rect 95663 18560 95669 18720
rect 94463 18520 95669 18560
rect 95721 18520 95727 18720
rect 94463 18397 94475 18520
rect 94399 18391 94475 18397
rect 94633 18424 95310 18438
rect 94414 18384 94454 18391
rect 94633 18387 95299 18424
rect 94633 18279 94684 18387
rect 93698 18228 94684 18279
rect 94789 18330 94853 18351
rect 92200 18129 92265 18130
rect 92201 18128 92265 18129
rect 94789 18130 94795 18330
rect 94847 18130 94853 18330
rect 95293 18264 95299 18387
rect 95287 18224 95299 18264
rect 95351 18224 95357 18424
rect 94789 18128 94853 18130
rect 88753 17913 93083 18072
rect 94358 17913 95047 18072
rect 88753 17899 95047 17913
rect 89235 17386 89245 17441
rect 89300 17386 95389 17441
rect 95444 17386 95453 17441
rect 89405 17305 89418 17357
rect 89470 17305 95561 17357
rect 89405 17302 95561 17305
rect 95616 17302 95623 17357
rect 89493 17271 95666 17273
rect 89493 17219 89503 17271
rect 89555 17219 95666 17271
rect 89493 17218 95666 17219
rect 95721 17218 95728 17273
rect 95933 17189 95969 23432
rect 96021 17189 96049 25402
rect 97096 25396 97150 25402
rect 96150 25192 96288 25239
rect 96150 21287 96194 25192
rect 96253 21287 96288 25192
rect 96150 19645 96166 21287
rect 96273 19645 96288 21287
rect 96150 17415 96194 19645
rect 96253 17415 96288 19645
rect 138094 25192 138232 25239
rect 138094 21287 138129 25192
rect 138188 21287 138232 25192
rect 138094 20345 138109 21287
rect 138216 20345 138232 21287
rect 138094 19955 138129 20345
rect 138188 19955 138232 20345
rect 138094 19645 138109 19955
rect 138216 19645 138232 19955
rect 96150 17364 96288 17415
rect 97102 17515 97150 17623
rect 97102 17463 97151 17515
rect 89574 17186 95174 17189
rect 89574 17134 89587 17186
rect 89639 17134 95174 17186
rect 95229 17134 95246 17189
rect 95933 17147 96049 17189
rect 89660 17103 95292 17105
rect 89660 17051 89671 17103
rect 89723 17051 95292 17103
rect 89660 17050 95292 17051
rect 95347 17050 95356 17105
rect 97102 17000 97150 17463
rect 91319 16872 91325 16926
rect 91379 16872 92207 16926
rect 92261 16872 92267 16926
rect 92466 16897 92472 16949
rect 92524 16947 92530 16949
rect 97097 16947 97150 17000
rect 92524 16899 97150 16947
rect 92524 16897 92530 16899
rect 92586 16801 92592 16853
rect 92644 16851 92650 16853
rect 99237 16851 99285 17623
rect 92644 16803 99285 16851
rect 92644 16801 92650 16803
rect 94654 16704 94660 16756
rect 94712 16754 94718 16756
rect 103505 16754 103559 17703
rect 138094 17415 138129 19645
rect 138188 17415 138232 19645
rect 138094 17364 138232 17415
rect 138333 17189 138361 25402
rect 138413 24634 138449 25430
rect 138413 24602 138541 24634
rect 138413 23432 138541 23463
rect 138413 17189 138449 23432
rect 138333 17147 138449 17189
rect 138678 22753 138878 22796
rect 94712 16706 103559 16754
rect 94712 16704 94718 16706
rect 89326 16569 89332 16621
rect 89384 16615 89390 16621
rect 94469 16615 94475 16621
rect 89384 16575 94475 16615
rect 89384 16569 89390 16575
rect 94469 16569 94475 16575
rect 94527 16615 94533 16621
rect 94527 16575 118579 16615
rect 94527 16569 94533 16575
rect 94789 16481 94853 16484
rect 92377 16465 92429 16471
rect 91319 16384 91325 16438
rect 91379 16384 91385 16438
rect 94789 16429 94795 16481
rect 94847 16429 94853 16481
rect 94905 16435 94911 16487
rect 94963 16481 94969 16487
rect 94963 16441 101500 16481
rect 94963 16435 94969 16441
rect 94789 16424 94841 16429
rect 92377 16407 92429 16413
rect 89524 16035 89640 16077
rect 89524 9792 89560 16035
rect 89432 9761 89560 9792
rect 89432 8590 89560 8622
rect 89524 7794 89560 8590
rect 89612 7822 89640 16035
rect 89741 15809 89879 15860
rect 89741 13579 89785 15809
rect 89844 13579 89879 15809
rect 90792 15549 91008 15560
rect 90792 15439 90874 15549
rect 90993 15439 91008 15549
rect 91325 15439 91379 16384
rect 92383 15600 92423 16407
rect 94506 16366 94841 16424
rect 94506 15598 94564 16366
rect 101460 15579 101500 16441
rect 118539 15514 118579 16575
rect 138332 16035 138448 16077
rect 138093 15809 138231 15860
rect 137230 15709 137302 15761
rect 90792 15424 91008 15439
rect 89741 11937 89757 13579
rect 89864 11937 89879 13579
rect 89741 8032 89785 11937
rect 89844 8032 89879 11937
rect 138093 13579 138128 15809
rect 138187 13579 138231 15809
rect 138093 13261 138108 13579
rect 138215 13261 138231 13579
rect 138093 12821 138128 13261
rect 138187 12821 138231 13261
rect 138093 11937 138108 12821
rect 138215 11937 138231 12821
rect 91043 8682 91095 8886
rect 90772 8630 91095 8682
rect 89741 7985 89879 8032
rect 138093 8032 138128 11937
rect 138187 8032 138231 11937
rect 138093 7985 138231 8032
rect 138332 7822 138360 16035
rect 138412 9792 138448 16035
rect 138678 10827 138878 22369
rect 138412 9761 138540 9792
rect 89612 7803 138360 7822
rect 89612 7794 89665 7803
rect 89524 7759 89665 7794
rect 138307 7794 138360 7803
rect 138412 8590 138540 8622
rect 138412 7794 138448 8590
rect 138307 7759 138448 7794
rect 89524 7744 138448 7759
rect 89241 7180 89247 7185
rect 89234 7137 89247 7180
rect 89241 7133 89247 7137
rect 89299 7180 89305 7185
rect 90409 7180 90415 7185
rect 89299 7137 90415 7180
rect 89299 7133 89305 7137
rect 90409 7133 90415 7137
rect 90467 7180 90473 7185
rect 90467 7137 90475 7180
rect 90467 7133 90473 7137
rect 89524 6978 138448 6993
rect 89524 6943 89665 6978
rect 89524 6147 89560 6943
rect 89432 6115 89560 6147
rect 89612 6934 89665 6943
rect 90370 6934 90560 6978
rect 138307 6943 138448 6978
rect 138307 6934 138360 6943
rect 89612 6915 138360 6934
rect 89432 4945 89560 4976
rect 89524 -1298 89560 4945
rect 89612 -1298 89640 6915
rect 89741 6705 89879 6752
rect 89741 2800 89785 6705
rect 89844 2800 89879 6705
rect 89741 1158 89757 2800
rect 89864 1158 89879 2800
rect 89741 -1072 89785 1158
rect 89844 -1072 89879 1158
rect 89741 -1123 89879 -1072
rect 138093 6705 138231 6752
rect 138093 2800 138128 6705
rect 138187 2800 138231 6705
rect 138093 1891 138108 2800
rect 138215 1891 138231 2800
rect 138093 1451 138128 1891
rect 138187 1451 138231 1891
rect 138093 1158 138108 1451
rect 138215 1158 138231 1451
rect 138093 -1072 138128 1158
rect 138187 -1072 138231 1158
rect 138093 -1123 138231 -1072
rect 89524 -1340 89640 -1298
rect 138332 -1298 138360 6915
rect 138412 6147 138448 6943
rect 138412 6115 138540 6147
rect 138412 4945 138540 4976
rect 138412 -1298 138448 4945
rect 138332 -1340 138448 -1298
rect 138678 4349 138878 10443
rect 89242 -1460 89248 -1408
rect 89300 -1415 89306 -1408
rect 89300 -1455 138018 -1415
rect 89300 -1460 89306 -1455
rect 137613 -9998 137619 -9946
rect 137671 -9952 137677 -9946
rect 137978 -9952 138018 -1455
rect 138332 -2445 138448 -2403
rect 137671 -9992 138018 -9952
rect 138093 -2671 138231 -2620
rect 138093 -4901 138128 -2671
rect 138187 -4901 138231 -2671
rect 138093 -5165 138108 -4901
rect 138215 -5165 138231 -4901
rect 138093 -5608 138128 -5165
rect 138187 -5608 138231 -5165
rect 138093 -6543 138108 -5608
rect 138215 -6543 138231 -5608
rect 137671 -9998 137677 -9992
rect 138093 -10448 138128 -6543
rect 138187 -10448 138231 -6543
rect 138093 -10495 138231 -10448
rect 138332 -10658 138360 -2445
rect 138412 -8688 138448 -2445
rect 138678 -7626 138878 3965
rect 138998 20373 139198 20427
rect 138998 13240 139198 19989
rect 138998 1870 139198 12856
rect 138998 -5249 139198 1486
rect 139318 19525 139518 19570
rect 139318 14153 139518 19141
rect 139318 1018 139518 13769
rect 139318 -4387 139518 634
rect 139318 -4812 139518 -4771
rect 138998 -5669 139198 -5633
rect 138678 -8051 138878 -8010
rect 138412 -8719 138540 -8688
rect 135144 -10677 138360 -10658
rect 135144 -10721 135416 -10677
rect 138307 -10686 138360 -10677
rect 138412 -9890 138540 -9858
rect 138412 -10686 138448 -9890
rect 138307 -10721 138448 -10686
rect 135144 -10736 138448 -10721
<< via1 >>
rect 93088 24381 94360 24496
rect 90131 24062 90264 24164
rect 92723 24062 92856 24164
rect 89122 23825 89505 23882
rect 90501 23564 91780 23781
rect 92696 23282 92748 23334
rect 92207 23204 92259 23214
rect 92207 23025 92252 23204
rect 92252 23025 92259 23204
rect 95391 23404 95443 23604
rect 95788 23463 95969 24602
rect 95969 23463 96002 24602
rect 92207 23014 92259 23025
rect 94795 23204 94847 23214
rect 94795 23025 94798 23204
rect 94798 23025 94844 23204
rect 94844 23025 94847 23204
rect 94795 23014 94847 23025
rect 95740 23127 95792 23327
rect 93083 22753 94353 22968
rect 90131 22434 90264 22536
rect 92723 22434 92856 22536
rect 89122 22197 89505 22254
rect 90501 21938 91780 22155
rect 92740 21671 92792 21723
rect 92207 21576 92259 21586
rect 92207 21397 92252 21576
rect 92252 21397 92259 21576
rect 95481 21776 95533 21976
rect 95719 21776 95771 21976
rect 94795 21576 94847 21586
rect 92207 21386 92259 21397
rect 94795 21397 94798 21576
rect 94798 21397 94844 21576
rect 94844 21397 94847 21576
rect 94795 21386 94847 21397
rect 95060 21493 95112 21693
rect 95593 21500 95645 21700
rect 93087 21120 94357 21335
rect 90131 20806 90264 20908
rect 92723 20806 92856 20908
rect 89125 20569 89505 20626
rect 90505 20307 91784 20524
rect 92730 20084 92782 20136
rect 95563 20148 95615 20348
rect 92207 19948 92259 19958
rect 92207 19769 92252 19948
rect 92252 19769 92259 19948
rect 92207 19758 92259 19769
rect 94795 19948 94847 19958
rect 94795 19769 94798 19948
rect 94798 19769 94844 19948
rect 94844 19769 94847 19948
rect 94795 19758 94847 19769
rect 95183 19856 95235 20056
rect 93085 19500 94355 19715
rect 90131 19178 90264 19280
rect 92723 19178 92856 19280
rect 89129 18941 89505 18998
rect 90501 18680 91780 18897
rect 92699 18433 92751 18485
rect 92207 18320 92259 18330
rect 92207 18141 92252 18320
rect 92252 18141 92259 18320
rect 92207 18130 92259 18141
rect 95669 18520 95721 18720
rect 94795 18320 94847 18330
rect 94795 18141 94798 18320
rect 94798 18141 94844 18320
rect 94844 18141 94847 18320
rect 94795 18130 94847 18141
rect 95299 18224 95351 18424
rect 93083 17913 94358 18076
rect 89245 17386 89300 17441
rect 95389 17386 95444 17441
rect 89418 17305 89470 17357
rect 95561 17302 95616 17357
rect 89503 17219 89555 17271
rect 95666 17218 95721 17273
rect 96166 19645 96194 21287
rect 96194 19645 96253 21287
rect 96253 19645 96273 21287
rect 138109 20345 138129 21287
rect 138129 20345 138188 21287
rect 138188 20345 138216 21287
rect 138109 19645 138129 19955
rect 138129 19645 138188 19955
rect 138188 19645 138216 19955
rect 89587 17134 89639 17186
rect 95174 17134 95229 17189
rect 89671 17051 89723 17103
rect 95292 17050 95347 17105
rect 91325 16872 91379 16926
rect 92207 16872 92261 16926
rect 92472 16897 92524 16949
rect 92592 16801 92644 16853
rect 94660 16704 94712 16756
rect 138380 23463 138413 24602
rect 138413 23463 138541 24602
rect 138678 22369 138878 22753
rect 89332 16569 89384 16621
rect 94475 16569 94527 16621
rect 91325 16384 91379 16438
rect 92377 16413 92429 16465
rect 94795 16429 94847 16481
rect 94911 16435 94963 16487
rect 89432 8622 89560 9761
rect 89560 8622 89593 9761
rect 89757 11937 89785 13579
rect 89785 11937 89844 13579
rect 89844 11937 89864 13579
rect 138108 13261 138128 13579
rect 138128 13261 138187 13579
rect 138187 13261 138215 13579
rect 138108 11937 138128 12821
rect 138128 11937 138187 12821
rect 138187 11937 138215 12821
rect 138678 10443 138878 10827
rect 138379 8622 138412 9761
rect 138412 8622 138540 9761
rect 89247 7133 89299 7185
rect 90415 7133 90467 7185
rect 89432 4976 89560 6115
rect 89560 4976 89593 6115
rect 89757 1158 89785 2800
rect 89785 1158 89844 2800
rect 89844 1158 89864 2800
rect 138108 1891 138128 2800
rect 138128 1891 138187 2800
rect 138187 1891 138215 2800
rect 138108 1158 138128 1451
rect 138128 1158 138187 1451
rect 138187 1158 138215 1451
rect 138379 4976 138412 6115
rect 138412 4976 138540 6115
rect 138678 3965 138878 4349
rect 89248 -1460 89300 -1408
rect 137619 -9998 137671 -9946
rect 138108 -5165 138128 -4901
rect 138128 -5165 138187 -4901
rect 138187 -5165 138215 -4901
rect 138108 -6543 138128 -5608
rect 138128 -6543 138187 -5608
rect 138187 -6543 138215 -5608
rect 138998 19989 139198 20373
rect 138998 12856 139198 13240
rect 138998 1486 139198 1870
rect 139318 19141 139518 19525
rect 139318 13769 139518 14153
rect 139318 634 139518 1018
rect 139318 -4771 139518 -4387
rect 138998 -5633 139198 -5249
rect 138678 -8010 138878 -7626
rect 138379 -9858 138412 -8719
rect 138412 -9858 138540 -8719
<< metal2 >>
rect 89111 23882 89505 24643
rect 89111 23825 89122 23882
rect 89111 22254 89505 23825
rect 89111 22197 89122 22254
rect 89111 20626 89505 22197
rect 89111 20569 89125 20626
rect 89111 19231 89505 20569
rect 89111 18998 89142 19231
rect 89474 18998 89505 19231
rect 89750 19245 89790 25266
rect 89870 20887 89910 25266
rect 89990 22510 90030 25266
rect 90110 24180 90150 25266
rect 90110 24164 90280 24180
rect 90110 24062 90131 24164
rect 90264 24062 90280 24164
rect 90110 24046 90280 24062
rect 90488 23781 91793 24554
rect 90488 23564 90501 23781
rect 91780 23564 91793 23781
rect 90110 22536 90280 22552
rect 90110 22510 90131 22536
rect 89990 22470 90131 22510
rect 90110 22434 90131 22470
rect 90264 22434 90280 22536
rect 90110 22418 90280 22434
rect 90488 22155 91793 23564
rect 92207 23214 92259 23222
rect 92207 23004 92259 23014
rect 90488 21938 90501 22155
rect 91780 21938 91793 22155
rect 90488 21255 91793 21938
rect 92213 21738 92253 23004
rect 92342 22218 92382 25266
rect 92462 22339 92502 25266
rect 92578 24848 92618 25266
rect 92578 22510 92622 24848
rect 92702 24180 92742 25266
rect 97246 24913 137385 25101
rect 97081 24760 98770 24845
rect 99241 24777 103040 24845
rect 99209 24773 103040 24777
rect 95606 24721 98770 24760
rect 93070 24604 94373 24644
rect 93070 24496 93104 24604
rect 94346 24496 94373 24604
rect 93070 24381 93088 24496
rect 94360 24381 94373 24496
rect 92702 24164 92872 24180
rect 92702 24062 92723 24164
rect 92856 24062 92872 24164
rect 92702 24046 92872 24062
rect 92702 23340 92742 24046
rect 93070 23459 93104 24381
rect 94346 23459 94373 24381
rect 95397 23610 95437 23632
rect 92696 23334 92748 23340
rect 92696 23276 92748 23282
rect 93070 22968 94373 23459
rect 95391 23604 95443 23610
rect 95391 23396 95443 23404
rect 94795 23214 94847 23222
rect 94795 23004 94847 23014
rect 93070 22753 93083 22968
rect 94353 22753 94373 22968
rect 92702 22536 92872 22552
rect 92702 22510 92723 22536
rect 92578 22470 92723 22510
rect 92702 22434 92723 22470
rect 92856 22434 92872 22536
rect 92702 22418 92872 22434
rect 92462 22299 92641 22339
rect 92342 22178 92522 22218
rect 92213 21698 92364 21738
rect 92207 21586 92259 21594
rect 92207 21376 92259 21386
rect 90110 20908 90280 20924
rect 90110 20887 90131 20908
rect 89870 20847 90131 20887
rect 90110 20806 90131 20847
rect 90264 20806 90280 20908
rect 90110 20790 90280 20806
rect 90488 20524 90532 21255
rect 91734 20524 91793 21255
rect 90488 20307 90505 20524
rect 91784 20307 91793 20524
rect 90488 19664 90532 20307
rect 91734 19664 91793 20307
rect 92213 20197 92253 21376
rect 92324 20543 92364 21698
rect 92482 20770 92522 22178
rect 92601 20887 92641 22299
rect 92746 21729 92786 22418
rect 92740 21723 92792 21729
rect 92740 21665 92792 21671
rect 93070 21335 94373 22753
rect 94801 21894 94841 23004
rect 93070 21120 93087 21335
rect 94357 21120 94373 21335
rect 92702 20908 92872 20924
rect 92702 20887 92723 20908
rect 92601 20847 92723 20887
rect 92702 20806 92723 20847
rect 92856 20806 92872 20908
rect 92702 20790 92872 20806
rect 92482 20730 92642 20770
rect 92324 20503 92493 20543
rect 92213 20157 92383 20197
rect 92207 19958 92259 19966
rect 92207 19748 92259 19758
rect 90110 19280 90280 19296
rect 90110 19245 90131 19280
rect 89750 19205 90131 19245
rect 90110 19178 90131 19205
rect 90264 19178 90280 19280
rect 90110 19162 90280 19178
rect 89111 18941 89129 18998
rect 89111 18093 89142 18941
rect 89474 18093 89505 18941
rect 89111 17850 89505 18093
rect 90488 18897 91793 19664
rect 90488 18680 90501 18897
rect 91780 18680 91793 18897
rect 92213 18790 92253 19748
rect 92343 18956 92383 20157
rect 92453 19109 92493 20503
rect 92602 19245 92642 20730
rect 92736 20142 92776 20790
rect 92730 20136 92782 20142
rect 92730 20078 92782 20084
rect 93070 19715 94373 21120
rect 93070 19500 93085 19715
rect 94355 19500 94373 19715
rect 92702 19280 92872 19296
rect 92702 19245 92723 19280
rect 92602 19205 92723 19245
rect 92702 19178 92723 19205
rect 92856 19178 92872 19280
rect 92702 19162 92872 19178
rect 92453 19069 92637 19109
rect 92343 18916 92518 18956
rect 92213 18750 92391 18790
rect 90488 17843 91793 18680
rect 92207 18330 92259 18338
rect 92207 18120 92259 18130
rect 89250 17447 89298 17450
rect 89245 17441 89300 17447
rect 89245 17380 89300 17386
rect 89250 8466 89298 17380
rect 89418 17357 89470 17363
rect 89418 17299 89470 17305
rect 89334 16627 89382 16631
rect 89332 16621 89384 16627
rect 89332 16563 89384 16569
rect 89244 8457 89300 8466
rect 89244 8392 89300 8401
rect 89250 7191 89298 8392
rect 89247 7185 89299 7191
rect 89247 7127 89299 7133
rect 89250 -1402 89298 7127
rect 89334 -745 89382 16563
rect 89418 10838 89469 17299
rect 89503 17271 89555 17277
rect 89503 17213 89555 17219
rect 89505 10922 89553 17213
rect 89587 17186 89639 17192
rect 89587 17128 89639 17134
rect 89589 11006 89637 17128
rect 89671 17103 89723 17109
rect 89671 17045 89723 17051
rect 89673 13808 89721 17045
rect 92213 16932 92253 18120
rect 91325 16926 91379 16932
rect 91325 16438 91379 16872
rect 92207 16926 92261 16932
rect 92207 16866 92261 16872
rect 92213 16862 92253 16866
rect 92351 16465 92391 18750
rect 92478 16955 92518 18916
rect 92472 16949 92524 16955
rect 92472 16891 92524 16897
rect 92478 16886 92518 16891
rect 92597 16859 92637 19069
rect 92705 18491 92745 19162
rect 92699 18485 92751 18491
rect 92699 18427 92751 18433
rect 93070 18076 94373 19500
rect 93070 17913 93083 18076
rect 94358 17913 94373 18076
rect 93070 17858 94373 17913
rect 94481 21854 94841 21894
rect 92592 16853 92644 16859
rect 92592 16795 92644 16801
rect 92597 16785 92637 16795
rect 94481 16627 94521 21854
rect 95058 21693 95116 21701
rect 94795 21586 94847 21594
rect 95058 21493 95060 21693
rect 95112 21493 95116 21693
rect 95058 21486 95117 21493
rect 94795 21376 94847 21386
rect 94801 20114 94841 21376
rect 94667 20074 94841 20114
rect 94667 16762 94707 20074
rect 94795 19958 94847 19966
rect 94795 19748 94847 19758
rect 94801 18806 94841 19748
rect 94801 18766 94957 18806
rect 94917 18600 94957 18766
rect 94917 18560 94979 18600
rect 94795 18330 94847 18338
rect 94795 18120 94847 18130
rect 94660 16756 94712 16762
rect 94660 16698 94712 16704
rect 94475 16621 94527 16627
rect 94475 16563 94527 16569
rect 94801 16487 94841 18120
rect 94917 16493 94957 18560
rect 95078 17387 95117 21486
rect 95184 20069 95223 20082
rect 95184 20062 95229 20069
rect 95183 20056 95235 20062
rect 95183 19848 95235 19856
rect 95184 17195 95223 19848
rect 95300 18437 95339 18456
rect 95300 18430 95345 18437
rect 95299 18424 95351 18430
rect 95299 18216 95351 18224
rect 95174 17189 95229 17195
rect 95174 17128 95229 17134
rect 95184 17127 95223 17128
rect 95300 17111 95339 18216
rect 95397 17447 95437 23396
rect 95606 23184 95646 24721
rect 97081 24657 98770 24721
rect 99058 24733 103040 24773
rect 95759 24602 96023 24634
rect 99058 24618 99098 24733
rect 99209 24657 103040 24733
rect 103322 24663 137385 24851
rect 95759 23463 95788 24602
rect 96002 23463 96023 24602
rect 95759 23432 96023 23463
rect 96239 24578 99098 24618
rect 95603 23124 95646 23184
rect 95740 23327 95792 23334
rect 96239 23311 96279 24578
rect 103322 24532 103362 24663
rect 95792 23271 96279 23311
rect 96345 24492 103362 24532
rect 138359 24602 138541 24634
rect 95481 21976 95533 21982
rect 95481 21768 95533 21776
rect 95487 17457 95527 21768
rect 95603 21740 95649 23124
rect 95740 23119 95792 23127
rect 96345 23005 96385 24492
rect 96784 24210 137661 24448
rect 138359 23463 138380 24602
rect 138359 23432 138541 23463
rect 95725 22965 96385 23005
rect 95725 21982 95765 22965
rect 138678 22753 138878 22777
rect 96784 22444 138678 22682
rect 138878 22444 138879 22682
rect 138678 22344 138878 22369
rect 95719 21976 95771 21982
rect 95719 21768 95771 21776
rect 95603 21709 95650 21740
rect 95591 21700 95650 21709
rect 95591 21500 95593 21700
rect 95645 21500 95649 21700
rect 126302 21567 137661 21702
rect 137335 21565 137661 21567
rect 95591 21493 95649 21500
rect 137413 21481 137661 21565
rect 126302 21464 137661 21481
rect 96111 21287 96302 21306
rect 95569 20354 95609 20378
rect 95563 20348 95615 20354
rect 95563 20140 95615 20148
rect 95389 17441 95444 17447
rect 95389 17380 95444 17386
rect 95397 17378 95437 17380
rect 95569 17363 95609 20140
rect 96111 19645 96166 21287
rect 96273 19645 96302 21287
rect 138080 21287 138271 21306
rect 96443 21022 96472 21256
rect 96727 21022 96773 21256
rect 137413 21172 137655 21256
rect 137545 21022 137655 21172
rect 137910 21022 137939 21256
rect 138080 20345 138109 21287
rect 138216 20345 138271 21287
rect 138998 20373 139198 20397
rect 96765 20076 138998 20310
rect 139198 20076 139201 20310
rect 138998 19964 139198 19989
rect 96111 19622 96302 19645
rect 138080 19645 138109 19955
rect 138216 19645 138271 19955
rect 138080 19622 138271 19645
rect 139318 19525 139518 19549
rect 137541 19411 139318 19412
rect 96765 19177 139318 19411
rect 139318 19116 139518 19141
rect 95675 18726 95715 18740
rect 95669 18720 95721 18726
rect 95669 18512 95721 18520
rect 95561 17357 95616 17363
rect 95561 17296 95616 17302
rect 95569 17294 95609 17296
rect 95675 17279 95715 18512
rect 96442 18284 96471 18518
rect 96726 18284 96773 18518
rect 137500 18284 137661 18518
rect 137911 18284 137940 18518
rect 96765 17949 137500 18187
rect 97092 17554 98763 17786
rect 99226 17554 103040 17786
rect 103482 17554 137257 17786
rect 97267 17284 137417 17479
rect 95666 17273 95721 17279
rect 97268 17247 137417 17284
rect 95666 17212 95721 17218
rect 95675 17211 95715 17212
rect 95292 17105 95347 17111
rect 95292 17044 95347 17050
rect 95300 17043 95339 17044
rect 94911 16487 94963 16493
rect 94795 16481 94847 16487
rect 92351 16419 92377 16465
rect 92371 16413 92377 16419
rect 92429 16413 92435 16465
rect 94911 16429 94963 16435
rect 94795 16423 94847 16429
rect 91325 16375 91379 16384
rect 90556 15746 137113 15977
rect 90556 15745 103128 15746
rect 90716 15438 90828 15670
rect 91270 15438 91374 15670
rect 91816 15438 92444 15670
rect 92860 15438 100992 15670
rect 101408 15438 118076 15670
rect 118504 15438 137292 15670
rect 90436 15271 137604 15275
rect 90436 15037 137610 15271
rect 90033 14706 90062 14940
rect 90317 14706 90436 14940
rect 137610 14706 137655 14940
rect 137910 14706 137939 14940
rect 139318 14153 139518 14177
rect 90312 13814 139318 14048
rect 90312 13813 90432 13814
rect 89673 13760 89996 13808
rect 89702 13579 89893 13602
rect 89702 11937 89757 13579
rect 89864 11937 89893 13579
rect 89702 11918 89893 11937
rect 89948 11790 89996 13760
rect 139518 13814 139522 14048
rect 139318 13744 139518 13769
rect 138079 13579 138270 13602
rect 138079 13261 138108 13579
rect 138215 13261 138270 13579
rect 138998 13240 139198 13264
rect 90356 12914 138998 13148
rect 138997 12856 138998 12914
rect 139198 12912 139208 13146
rect 138997 12854 139198 12856
rect 138998 12831 139198 12854
rect 90034 11968 90063 12202
rect 90318 12068 90432 12202
rect 90441 12068 90560 12078
rect 90318 11994 90560 12068
rect 90318 11984 90441 11994
rect 90318 11968 90432 11984
rect 137608 11968 137654 12202
rect 137909 11968 137938 12202
rect 138079 11937 138108 12821
rect 138215 11937 138270 12821
rect 138079 11918 138270 11937
rect 89916 11742 89996 11790
rect 90312 11743 108079 11760
rect 89589 10958 89880 11006
rect 89505 10874 89796 10922
rect 89418 10788 89712 10838
rect 89432 9761 89614 9792
rect 89593 8622 89614 9761
rect 89432 8590 89614 8622
rect 89664 8338 89712 10788
rect 89658 8329 89718 8338
rect 89658 8260 89718 8269
rect 89748 8198 89796 10874
rect 89742 8189 89802 8198
rect 89742 8120 89802 8129
rect 89832 8069 89880 10958
rect 89826 8060 89886 8069
rect 89826 7991 89886 8000
rect 89916 7939 89964 11742
rect 90312 11659 90560 11743
rect 90312 11657 90638 11659
rect 90312 11522 108079 11657
rect 138678 10827 138878 10851
rect 90368 10543 138678 10781
rect 138878 10498 138879 10736
rect 138678 10418 138878 10443
rect 138358 9761 138540 9792
rect 90312 8776 137597 9014
rect 138358 8622 138379 9761
rect 138358 8590 138540 8622
rect 91272 8478 91392 8567
rect 91272 8422 91306 8478
rect 91362 8422 91392 8478
rect 91272 8379 91392 8422
rect 91818 8491 92456 8567
rect 91818 8435 91846 8491
rect 91902 8435 92456 8491
rect 91818 8379 92456 8435
rect 92882 8491 100978 8567
rect 92882 8435 92911 8491
rect 92967 8435 100978 8491
rect 92882 8379 100978 8435
rect 101400 8495 118082 8567
rect 101400 8439 101452 8495
rect 101508 8439 118082 8495
rect 101400 8379 118082 8439
rect 118510 8494 137300 8567
rect 118510 8438 118542 8494
rect 118598 8438 137300 8494
rect 118510 8379 137300 8438
rect 90751 8311 90846 8317
rect 90588 8123 137135 8311
rect 89910 7930 89970 7939
rect 89910 7861 89970 7870
rect 90415 7185 90467 7191
rect 90415 7127 90467 7133
rect 90420 6338 90463 7127
rect 90588 6426 137135 6614
rect 90751 6338 137300 6358
rect 90420 6295 137300 6338
rect 90751 6170 137300 6295
rect 89432 6115 89614 6147
rect 89593 4976 89614 6115
rect 138358 6115 138540 6147
rect 90312 5723 137597 5961
rect 89432 4945 89614 4976
rect 138358 4976 138379 6115
rect 138358 4945 138540 4976
rect 138678 4349 138878 4373
rect 90368 3965 138678 4194
rect 138878 4001 138879 4239
rect 90368 3956 138878 3965
rect 138678 3940 138878 3956
rect 90312 3080 108079 3215
rect 90312 3078 90638 3080
rect 90312 2994 90560 3078
rect 90312 2977 108079 2994
rect 89702 2800 89893 2819
rect 89702 1158 89757 2800
rect 89864 1158 89893 2800
rect 90034 2585 90063 2819
rect 90318 2803 90364 2819
rect 90318 2719 90560 2803
rect 138079 2800 138270 2819
rect 90318 2585 90364 2719
rect 137608 2535 137654 2769
rect 137909 2535 137938 2769
rect 138079 1891 138108 2800
rect 138215 1891 138270 2800
rect 138998 1870 139198 1894
rect 90356 1589 138998 1823
rect 139198 1531 139204 1765
rect 138998 1461 139198 1486
rect 89702 1135 89893 1158
rect 138079 1158 138108 1451
rect 138215 1158 138270 1451
rect 138079 1135 138270 1158
rect 139318 1018 139518 1042
rect 90312 924 90432 925
rect 90312 690 139318 924
rect 139318 609 139518 634
rect 90033 -203 90062 31
rect 90317 -203 90434 31
rect 137610 -203 137655 31
rect 137910 -203 137939 31
rect 90312 -538 137616 -300
rect 90716 -745 137845 -701
rect 89334 -793 137845 -745
rect 90716 -933 137845 -793
rect 90556 -1240 137113 -1008
rect 137789 -1114 137845 -933
rect 89248 -1408 89300 -1402
rect 89248 -1466 89300 -1460
rect 135412 -2735 137704 -2503
rect 137789 -2807 137846 -1114
rect 137624 -2810 137846 -2807
rect 135572 -2864 137846 -2810
rect 135572 -3042 137704 -2864
rect 135168 -3443 137704 -3205
rect 135168 -3774 135290 -3540
rect 137608 -3774 137655 -3540
rect 137910 -3774 137939 -3540
rect 139318 -4387 139518 -4363
rect 135168 -4667 139318 -4433
rect 139318 -4796 139518 -4771
rect 138079 -4901 138270 -4878
rect 138079 -5165 138108 -4901
rect 138215 -5165 138270 -4901
rect 138998 -5249 139198 -5225
rect 135224 -5566 138998 -5332
rect 137607 -6328 137654 -6278
rect 135214 -6462 137654 -6328
rect 135214 -6546 135416 -6462
rect 137392 -6512 137654 -6462
rect 137909 -6512 137938 -6278
rect 137392 -6546 137607 -6512
rect 135214 -6562 137607 -6546
rect 138079 -6543 138108 -5608
rect 138215 -6543 138270 -5608
rect 138998 -5658 139198 -5633
rect 138079 -6562 138270 -6543
rect 135168 -6737 137704 -6720
rect 135168 -6821 135416 -6737
rect 135168 -6823 135494 -6821
rect 137392 -6823 137704 -6737
rect 135168 -6958 137704 -6823
rect 138678 -7603 138878 -7602
rect 138677 -7626 138878 -7603
rect 138677 -7699 138678 -7626
rect 135224 -7937 138678 -7699
rect 138677 -8010 138678 -7937
rect 138878 -7937 138880 -7699
rect 138677 -8035 138878 -8010
rect 138358 -8719 138540 -8688
rect 135168 -9704 137704 -9466
rect 138358 -9858 138379 -8719
rect 138358 -9890 138540 -9858
rect 135607 -9946 137704 -9913
rect 135607 -9998 137619 -9946
rect 137671 -9998 137704 -9946
rect 135607 -10101 137704 -9998
rect 135444 -10357 137704 -10169
<< via2 >>
rect 89142 18998 89474 19231
rect 93104 24496 94346 24604
rect 93104 24381 94346 24496
rect 93104 23459 94346 24381
rect 90532 20524 91734 21255
rect 90532 20307 91734 20524
rect 90532 19664 91734 20307
rect 89142 18941 89474 18998
rect 89142 18093 89474 18941
rect 89244 8401 89300 8457
rect 95788 23463 96002 24602
rect 138380 23463 138541 24602
rect 125319 21565 137335 21567
rect 97234 21481 137413 21565
rect 96166 19645 96273 21287
rect 96472 21022 96727 21256
rect 97235 21156 137413 21240
rect 137655 21022 137910 21256
rect 138109 20345 138216 21287
rect 138109 19645 138216 19955
rect 96471 18284 96726 18518
rect 137661 18284 137911 18518
rect 90062 14706 90317 14940
rect 137655 14706 137910 14940
rect 89757 11937 89864 13579
rect 138108 13261 138215 13579
rect 90063 11968 90318 12202
rect 90560 11994 137146 12078
rect 137654 11968 137909 12202
rect 138108 11937 138215 12821
rect 89432 8622 89593 9761
rect 89658 8269 89718 8329
rect 89742 8129 89802 8189
rect 89826 8000 89886 8060
rect 90560 11659 137147 11743
rect 90638 11657 109062 11659
rect 138379 8622 138540 9761
rect 91306 8422 91362 8478
rect 91846 8435 91902 8491
rect 92911 8435 92967 8491
rect 101452 8439 101508 8495
rect 118542 8438 118598 8494
rect 89910 7870 89970 7930
rect 89432 4976 89593 6115
rect 138379 4976 138540 6115
rect 90638 3078 109062 3080
rect 90560 2994 137147 3078
rect 89757 1158 89864 2800
rect 90063 2585 90318 2819
rect 90560 2669 137146 2753
rect 137654 2535 137909 2769
rect 138108 1891 138215 2800
rect 138108 1158 138215 1451
rect 90062 -203 90317 31
rect 137655 -203 137910 31
rect 137655 -3774 137910 -3540
rect 138108 -5165 138215 -4901
rect 135416 -6546 137392 -6462
rect 137654 -6512 137909 -6278
rect 138108 -6543 138215 -5608
rect 135416 -6821 137392 -6737
rect 135494 -6823 137392 -6821
rect 138379 -9858 138540 -8719
<< metal3 >>
rect 93072 24604 94372 24631
rect 93072 23459 93104 24604
rect 94346 23459 94372 24604
rect 93072 23431 94372 23459
rect 95759 24602 96023 24634
rect 95759 23463 95788 24602
rect 96002 23463 96023 24602
rect 95759 23432 96023 23463
rect 90487 21255 91793 21308
rect 96461 21306 96739 24690
rect 138359 24602 138547 24634
rect 96842 21656 137538 21702
rect 96842 21654 125319 21656
rect 137335 21654 137538 21656
rect 96842 21480 97234 21654
rect 137413 21480 137538 21654
rect 96842 21464 137538 21480
rect 137643 21306 137921 24449
rect 138359 23463 138380 24602
rect 138541 23463 138547 24602
rect 138359 23432 138547 23463
rect 90487 19664 90532 21255
rect 91734 19664 91793 21255
rect 90487 19621 91793 19664
rect 96133 21287 96302 21306
rect 96133 19645 96166 21287
rect 96273 19645 96302 21287
rect 96133 19623 96302 19645
rect 96461 21291 137921 21306
rect 96461 21256 97234 21291
rect 96461 21022 96472 21256
rect 96727 21117 97234 21256
rect 137413 21256 137921 21291
rect 137413 21117 137655 21256
rect 96727 21072 137655 21117
rect 96727 21022 96739 21072
rect 89112 19231 89505 19260
rect 89112 18093 89142 19231
rect 89474 18093 89505 19231
rect 96461 18518 96739 21022
rect 96461 18284 96471 18518
rect 96726 18284 96739 18518
rect 96461 18247 96739 18284
rect 137643 21022 137655 21072
rect 137910 21022 137921 21256
rect 137643 18518 137921 21022
rect 138080 21287 138249 21306
rect 138080 19645 138109 21287
rect 138216 19645 138249 21287
rect 138080 19623 138249 19645
rect 137643 18284 137661 18518
rect 137911 18284 137921 18518
rect 137643 18251 137921 18284
rect 89112 18058 89505 18093
rect 90052 14940 90330 14977
rect 90052 14706 90062 14940
rect 90317 14706 90330 14940
rect 89724 13579 89893 13601
rect 89724 11937 89757 13579
rect 89864 11937 89893 13579
rect 89724 11918 89893 11937
rect 90052 12202 90330 14706
rect 90052 11968 90063 12202
rect 90318 12152 90330 12202
rect 137642 14940 137920 14977
rect 137642 14706 137655 14940
rect 137910 14706 137920 14940
rect 137642 12202 137920 14706
rect 137642 12152 137654 12202
rect 90318 12107 137654 12152
rect 90318 11968 90560 12107
rect 90052 11933 90560 11968
rect 137147 11968 137654 12107
rect 137909 11968 137920 12202
rect 137147 11933 137920 11968
rect 90052 11918 137920 11933
rect 138079 13579 138248 13601
rect 138079 11937 138108 13579
rect 138215 11937 138248 13579
rect 138079 11918 138248 11937
rect 89427 9761 89614 9792
rect 89427 8622 89432 9761
rect 89593 8622 89614 9761
rect 90052 8776 90330 11918
rect 90406 11744 137539 11760
rect 90406 11570 90560 11744
rect 137147 11570 137539 11744
rect 90406 11568 90638 11570
rect 109062 11568 137539 11570
rect 90406 11522 137539 11568
rect 90404 8930 93370 8990
rect 89427 8590 89614 8622
rect 89239 8459 89305 8462
rect 90404 8459 90464 8930
rect 89239 8457 90464 8459
rect 89239 8401 89244 8457
rect 89300 8401 90464 8457
rect 89239 8399 90464 8401
rect 90524 8810 93209 8870
rect 89239 8396 89305 8399
rect 89653 8329 89723 8334
rect 90524 8329 90584 8810
rect 89651 8269 89658 8329
rect 89718 8269 90584 8329
rect 90644 8670 92638 8730
rect 89653 8264 89723 8269
rect 89737 8189 89807 8194
rect 90644 8189 90704 8670
rect 89736 8129 89742 8189
rect 89802 8129 90704 8189
rect 90764 8550 91540 8610
rect 89737 8124 89807 8129
rect 89821 8060 89891 8065
rect 89821 8059 89826 8060
rect 89815 8000 89826 8059
rect 89886 8059 89891 8060
rect 90764 8059 90824 8550
rect 91480 8493 91540 8550
rect 91841 8493 91907 8496
rect 92578 8493 92638 8670
rect 93149 8497 93209 8810
rect 93310 8622 93370 8930
rect 137642 8774 137920 11918
rect 138358 9761 138545 9792
rect 138358 8622 138379 9761
rect 138540 8622 138545 9761
rect 93310 8562 101757 8622
rect 138358 8590 138545 8622
rect 101447 8497 101513 8500
rect 92906 8493 92972 8496
rect 91480 8491 91919 8493
rect 91301 8480 91367 8483
rect 89886 8000 90824 8059
rect 89815 7999 90824 8000
rect 90884 8478 91395 8480
rect 90884 8422 91306 8478
rect 91362 8422 91395 8478
rect 91480 8435 91846 8491
rect 91902 8435 91919 8491
rect 91480 8433 91919 8435
rect 92578 8491 92972 8493
rect 92578 8435 92911 8491
rect 92967 8435 92972 8491
rect 93149 8495 101516 8497
rect 93149 8439 101452 8495
rect 101508 8439 101516 8495
rect 93149 8437 101516 8439
rect 101697 8496 101757 8562
rect 118537 8496 118603 8499
rect 101697 8494 118608 8496
rect 101697 8438 118542 8494
rect 118598 8438 118608 8494
rect 92578 8433 92972 8435
rect 101447 8434 101513 8437
rect 101697 8436 118608 8438
rect 118537 8433 118603 8436
rect 91841 8430 91907 8433
rect 92906 8430 92972 8433
rect 90884 8420 91395 8422
rect 89821 7995 89891 7999
rect 89905 7930 89975 7935
rect 89905 7929 89910 7930
rect 89903 7870 89910 7929
rect 89970 7929 89975 7930
rect 90884 7929 90944 8420
rect 91301 8417 91367 8420
rect 89970 7870 90944 7929
rect 89903 7869 90944 7870
rect 89905 7865 89975 7869
rect 89427 6115 89614 6147
rect 89427 4976 89432 6115
rect 89593 4976 89614 6115
rect 89427 4945 89614 4976
rect 90052 2819 90330 6203
rect 138358 6115 138545 6147
rect 90417 3169 137539 3215
rect 90417 3167 90638 3169
rect 109062 3167 137539 3169
rect 90417 2993 90560 3167
rect 137147 2993 137539 3167
rect 90417 2977 137539 2993
rect 137642 2819 137920 5968
rect 138358 4976 138379 6115
rect 138540 4976 138545 6115
rect 138358 4945 138545 4976
rect 89724 2800 89893 2819
rect 89724 1158 89757 2800
rect 89864 1158 89893 2800
rect 89724 1136 89893 1158
rect 90052 2585 90063 2819
rect 90318 2804 137920 2819
rect 90318 2630 90560 2804
rect 137147 2769 137920 2804
rect 137147 2630 137654 2769
rect 90318 2585 137654 2630
rect 90052 31 90330 2585
rect 90052 -203 90062 31
rect 90317 -203 90330 31
rect 90052 -240 90330 -203
rect 137642 2535 137654 2585
rect 137909 2535 137920 2769
rect 137642 31 137920 2535
rect 138079 2800 138248 2819
rect 138079 1158 138108 2800
rect 138215 1158 138248 2800
rect 138079 1136 138248 1158
rect 137642 -203 137655 31
rect 137910 -203 137920 31
rect 137642 -240 137920 -203
rect 137642 -3540 137920 -3503
rect 137642 -3774 137655 -3540
rect 137910 -3774 137920 -3540
rect 137642 -6278 137920 -3774
rect 135208 -6373 137516 -6328
rect 135208 -6547 135416 -6373
rect 137392 -6547 137516 -6373
rect 135208 -6562 137516 -6547
rect 137642 -6512 137654 -6278
rect 137909 -6512 137920 -6278
rect 135219 -6736 137516 -6720
rect 135219 -6910 135416 -6736
rect 135219 -6912 135494 -6910
rect 137392 -6912 137516 -6736
rect 135219 -6958 137516 -6912
rect 137642 -9703 137920 -6512
rect 138079 -4901 138248 -4879
rect 138079 -6543 138108 -4901
rect 138215 -6543 138248 -4901
rect 138079 -6562 138248 -6543
rect 138358 -8719 138545 -8688
rect 138358 -9858 138379 -8719
rect 138540 -9858 138545 -8719
rect 138358 -9890 138545 -9858
<< via3 >>
rect 93104 23459 94346 24604
rect 95788 23463 96002 24602
rect 125319 21654 137335 21656
rect 97234 21567 137413 21654
rect 97234 21565 125319 21567
rect 125319 21565 137335 21567
rect 137335 21565 137413 21567
rect 97234 21481 137413 21565
rect 97234 21480 137413 21481
rect 138380 23463 138541 24602
rect 90532 19664 91734 21255
rect 96166 19645 96273 21287
rect 97234 21240 137413 21291
rect 97234 21156 97235 21240
rect 97235 21156 137413 21240
rect 97234 21117 137413 21156
rect 89150 18093 89474 19231
rect 138109 20345 138216 21287
rect 138109 19955 138216 20345
rect 138109 19645 138216 19955
rect 89757 11937 89864 13579
rect 90560 12078 137147 12107
rect 90560 11994 137146 12078
rect 137146 11994 137147 12078
rect 90560 11933 137147 11994
rect 138108 13261 138215 13579
rect 138108 12821 138215 13261
rect 138108 11937 138215 12821
rect 89432 8622 89593 9761
rect 90560 11743 137147 11744
rect 90560 11659 137147 11743
rect 90560 11657 90638 11659
rect 90638 11657 109062 11659
rect 109062 11657 137147 11659
rect 90560 11570 137147 11657
rect 90638 11568 109062 11570
rect 138379 8622 138540 9761
rect 89432 4976 89593 6115
rect 90638 3167 109062 3169
rect 90560 3080 137147 3167
rect 90560 3078 90638 3080
rect 90638 3078 109062 3080
rect 109062 3078 137147 3080
rect 90560 2994 137147 3078
rect 90560 2993 137147 2994
rect 138379 4976 138540 6115
rect 89757 1158 89864 2800
rect 90560 2753 137147 2804
rect 90560 2669 137146 2753
rect 137146 2669 137147 2753
rect 90560 2630 137147 2669
rect 138108 1891 138215 2800
rect 138108 1451 138215 1891
rect 138108 1158 138215 1451
rect 135416 -6462 137392 -6373
rect 135416 -6546 137392 -6462
rect 135416 -6547 137392 -6546
rect 135416 -6737 137392 -6736
rect 135416 -6821 137392 -6737
rect 135416 -6823 135494 -6821
rect 135494 -6823 137392 -6821
rect 135416 -6910 137392 -6823
rect 135494 -6912 137392 -6910
rect 138108 -5165 138215 -4901
rect 138108 -5608 138215 -5165
rect 138108 -6543 138215 -5608
rect 138379 -9858 138540 -8719
<< metal4 >>
rect 88536 24604 96025 24633
rect 88536 23459 93104 24604
rect 94346 24602 96025 24604
rect 94346 23463 95788 24602
rect 96002 23463 96025 24602
rect 94346 23459 96025 23463
rect 88536 23433 96025 23459
rect 138357 24602 138545 24633
rect 138357 23463 138380 24602
rect 138541 23463 138545 24602
rect 138357 23433 138545 23463
rect 88536 21656 138541 23145
rect 88536 21654 125319 21656
rect 137335 21654 138541 21656
rect 88536 21480 97234 21654
rect 137413 21480 138541 21654
rect 88536 21460 138541 21480
rect 88536 21291 138541 21309
rect 88536 21287 97234 21291
rect 88536 21255 96166 21287
rect 88536 19664 90532 21255
rect 91734 19664 96166 21255
rect 88536 19645 96166 19664
rect 96273 21117 97234 21287
rect 137413 21287 138541 21291
rect 137413 21117 138109 21287
rect 96273 19645 138109 21117
rect 138216 19645 138541 21287
rect 88536 19624 138541 19645
rect 88536 19231 96025 19261
rect 88536 18093 89150 19231
rect 89474 18093 96025 19231
rect 88536 18061 96025 18093
rect 89432 13963 89616 15163
rect 89432 13579 138540 13600
rect 89432 11937 89757 13579
rect 89864 12107 138108 13579
rect 89864 11937 90560 12107
rect 89432 11933 90560 11937
rect 137147 11937 138108 12107
rect 138215 11937 138540 13579
rect 137147 11933 138540 11937
rect 89432 11915 138540 11933
rect 89432 11744 138540 11764
rect 89432 11570 90560 11744
rect 137147 11570 138540 11744
rect 89432 11568 90638 11570
rect 109062 11568 138540 11570
rect 89432 10079 138540 11568
rect 89429 9761 89616 9791
rect 89429 8622 89432 9761
rect 89593 8622 89616 9761
rect 89429 8591 89616 8622
rect 138356 9761 138544 9791
rect 138356 8622 138379 9761
rect 138540 8622 138544 9761
rect 138356 8591 138544 8622
rect 89429 6115 89616 6146
rect 89429 4976 89432 6115
rect 89593 4976 89616 6115
rect 89429 4946 89616 4976
rect 138356 6115 138543 6146
rect 138356 4976 138379 6115
rect 138540 4976 138543 6115
rect 138356 4946 138543 4976
rect 89432 3169 138540 4658
rect 89432 3167 90638 3169
rect 109062 3167 138540 3169
rect 89432 2993 90560 3167
rect 137147 2993 138540 3167
rect 89432 2973 138540 2993
rect 89432 2804 138540 2822
rect 89432 2800 90560 2804
rect 89432 1158 89757 2800
rect 89864 2630 90560 2800
rect 137147 2800 138540 2804
rect 137147 2630 138108 2800
rect 89864 1158 138108 2630
rect 138215 1158 138540 2800
rect 89432 1137 138540 1158
rect 89432 -426 89616 774
rect 135167 -4901 138540 -4880
rect 135167 -6373 138108 -4901
rect 135167 -6547 135416 -6373
rect 137392 -6543 138108 -6373
rect 138215 -6543 138540 -4901
rect 137392 -6547 138540 -6543
rect 135167 -6565 138540 -6547
rect 135168 -6736 138540 -6716
rect 135168 -6910 135416 -6736
rect 135168 -6912 135494 -6910
rect 137392 -6912 138540 -6736
rect 135168 -8401 138540 -6912
rect 138356 -8719 138546 -8689
rect 138356 -9858 138379 -8719
rect 138540 -9858 138546 -8719
rect 138356 -9889 138546 -9858
use bias_nstack  bias_nstack_0
array 0 75 -534 0 0 -4355
timestamp 1747745286
transform 1 0 133578 0 1 24324
box 3258 -2860 3926 785
use bias_nstack  bias_nstack_1
array 0 87 -534 0 0 -4355
timestamp 1747745286
transform -1 0 94395 0 -1 8900
box 3258 -2860 3926 785
use bias_nstack  bias_nstack_2
array 0 87 -534 0 0 -4355
timestamp 1747745286
transform -1 0 94395 0 1 5837
box 3258 -2860 3926 785
use bias_nstack  bias_nstack_3
array 0 3 -534 0 0 -4355
timestamp 1747745286
transform -1 0 139251 0 -1 -9580
box 3258 -2860 3926 785
use bias_pstack  bias_pstack_0
array 0 75 534 0 0 -4355
timestamp 1747752771
transform -1 0 139531 0 1 20918
box 1986 -3697 2714 338
use bias_pstack  bias_pstack_1
array 0 87 534 0 0 -4355
timestamp 1747752771
transform 1 0 88442 0 -1 12306
box 1986 -3697 2714 338
use bias_pstack  bias_pstack_2
array 0 87 534 0 0 -4355
timestamp 1747752771
transform 1 0 88442 0 1 2431
box 1986 -3697 2714 338
use bias_pstack  bias_pstack_3
array 0 3 534 0 0 -4355
timestamp 1747752771
transform 1 0 133298 0 -1 -6174
box 1986 -3697 2714 338
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_8 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1746753973
transform 1 0 91893 0 -1 24486
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_9
timestamp 1746753973
transform 1 0 91893 0 -1 21230
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_10
timestamp 1746753973
transform 1 0 91893 0 -1 22858
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_11
timestamp 1746753973
transform 1 0 94485 0 -1 24486
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_12
timestamp 1746753973
transform 1 0 91893 0 -1 19602
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_13
timestamp 1746753973
transform 1 0 94485 0 -1 19602
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_16
timestamp 1746753973
transform 1 0 94485 0 -1 21230
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_17
timestamp 1746753973
transform 1 0 94485 0 -1 22858
box -66 -43 450 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1746753973
transform 1 0 89589 0 -1 24486
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_1
timestamp 1746753973
transform 1 0 89589 0 1 22858
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_2
timestamp 1746753973
transform 1 0 89589 0 -1 19602
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_3
timestamp 1746753973
transform 1 0 89589 0 1 17974
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_4
timestamp 1746753973
transform 1 0 89589 0 -1 21230
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_5
timestamp 1746753973
transform 1 0 89589 0 1 19602
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_6
timestamp 1746753973
transform 1 0 89589 0 -1 22858
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_7
timestamp 1746753973
transform 1 0 89589 0 1 21230
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_8 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1746753973
transform 1 0 92277 0 -1 24486
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_9
timestamp 1746753973
transform 1 0 92277 0 -1 21230
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_10
timestamp 1746753973
transform 1 0 92277 0 -1 22858
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_11
timestamp 1746753973
transform 1 0 94869 0 -1 24486
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_12
timestamp 1746753973
transform 1 0 92277 0 -1 19602
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_13
timestamp 1746753973
transform 1 0 94869 0 -1 19602
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_16
timestamp 1746753973
transform 1 0 94869 0 -1 21230
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_17
timestamp 1746753973
transform 1 0 94869 0 -1 22858
box -66 -43 162 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1746753973
transform 1 0 94485 0 1 22858
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_1
timestamp 1746753973
transform 1 0 91893 0 1 22858
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_2
timestamp 1746753973
transform 1 0 94485 0 1 21230
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_3
timestamp 1746753973
transform 1 0 94485 0 1 19602
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_4
timestamp 1746753973
transform 1 0 91893 0 1 17974
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_7
timestamp 1746753973
transform 1 0 91893 0 1 21230
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_10
timestamp 1746753973
transform 1 0 94485 0 1 17974
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_11
timestamp 1746753973
transform 1 0 91893 0 1 19602
box -66 -43 546 897
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
array 0 1 -2592 0 3 1628
timestamp 1746753973
transform 1 0 92373 0 -1 24486
box -66 -43 2178 1671
<< labels >>
flabel metal4 90311 1137 90544 2822 0 FreeSans 1600 270 0 0 avdd
port 1 nsew
flabel metal4 90312 2973 90545 4658 0 FreeSans 1600 270 0 0 avss
port 2 nsew
flabel metal4 90311 11915 90544 13600 0 FreeSans 1600 90 0 0 avdd
port 1 nsew
flabel metal4 90312 10079 90545 11764 0 FreeSans 1600 90 0 0 avss
port 2 nsew
flabel metal4 137603 19624 137662 21309 0 FreeSans 1600 270 0 0 avdd
port 1 nsew
flabel metal4 137603 21460 137661 23145 0 FreeSans 1600 270 0 0 avss
port 2 nsew
flabel metal2 89750 24891 89790 25266 0 FreeSans 400 270 0 0 ena[0]
port 22 nsew
flabel metal2 89870 24891 89910 25266 0 FreeSans 400 270 0 0 ena[1]
port 23 nsew
flabel metal2 89990 24891 90030 25266 0 FreeSans 400 270 0 0 ena[2]
port 21 nsew
flabel metal2 90110 24891 90150 25266 0 FreeSans 400 270 0 0 ena[3]
port 20 nsew
flabel metal2 92342 24891 92382 25266 0 FreeSans 400 270 0 0 ena[4]
port 25 nsew
flabel metal2 92462 24891 92502 25266 0 FreeSans 400 270 0 0 ena[5]
port 24 nsew
flabel metal2 92578 24891 92618 25266 0 FreeSans 400 270 0 0 ena[6]
port 16 nsew
flabel metal2 92702 24866 92742 25266 0 FreeSans 400 270 0 0 ena[7]
port 26 nsew
flabel comment s 95318 17560 95318 17560 0 FreeSans 320 90 0 0 ena_bit0
flabel comment s 92230 17318 92230 17318 0 FreeSans 320 90 0 0 enb_bit0
flabel comment s 95206 17570 95206 17570 0 FreeSans 320 90 0 0 ena_bit1
flabel comment s 92366 17326 92366 17326 0 FreeSans 320 90 0 0 enb_bit1
flabel metal2 95100 17558 95100 17558 0 FreeSans 320 90 0 0 ena_bit2
flabel metal2 95690 17560 95690 17560 0 FreeSans 320 90 0 0 ena_bit4
flabel metal2 95588 17560 95588 17560 0 FreeSans 320 90 0 0 ena_bit5
flabel metal2 95514 17568 95514 17568 0 FreeSans 320 90 0 0 ena_bit6
flabel metal2 95412 17560 95412 17560 0 FreeSans 320 90 0 0 ena_bit7
flabel metal2 92496 17318 92496 17318 0 FreeSans 320 90 0 0 enb_bit2
flabel metal2 92616 17292 92616 17292 0 FreeSans 320 90 0 0 enb_bit3
flabel metal2 94830 17314 94830 17314 0 FreeSans 320 90 0 0 enb_bit4
flabel metal2 94942 17310 94942 17310 0 FreeSans 320 90 0 0 enb_bit5
flabel metal2 94692 17284 94692 17284 0 FreeSans 320 90 0 0 enb_bit6
flabel metal2 94494 17262 94494 17262 0 FreeSans 320 90 0 0 enb_bit7
flabel metal2 96249 24061 96249 24061 0 FreeSans 320 90 0 0 ena_bit3
flabel metal4 135167 -6565 135400 -4880 0 FreeSans 1600 90 0 0 avdd
port 1 nsew
flabel metal4 135168 -8401 135401 -6716 0 FreeSans 1600 90 0 0 avss
port 2 nsew
flabel metal4 88536 18061 89136 19261 0 FreeSans 3200 270 0 0 dvdd
port 3 nsew
flabel metal4 88536 19624 89136 21309 0 FreeSans 3200 270 0 0 avdd
port 1 nsew
flabel metal4 88536 21460 89136 23145 0 FreeSans 3200 270 0 0 avss
port 2 nsew
flabel metal4 88536 23433 89136 24633 0 FreeSans 3200 270 0 0 dvss
port 4 nsew
<< properties >>
string MASKHINTS_HVI 88550 17750 95280 17980 88550 24480 95280 24705 94835 17735 95280 24695
<< end >>
