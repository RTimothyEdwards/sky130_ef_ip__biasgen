** sch_path: /home/tim/gits/sky130_ef_ip__biasgen/xschem/bias_generator.sch
**.subckt bias_generator avdd ena ena_snk_2000 vbg ena_src_50 ena_snk_3700 ena_src_100 ena_snk_5000_2 src_200_0 ena_src_200_2
*+ src_10000_0 src_400 src_600 src_test0 src_test1 src_10000_1 src_100 src_200_2 src_50 src_200_1 ena_snk_5000_1 ena_src_200_1 ena_snk_5000_0
*+ snk_test1 snk_5000_2 snk_5000_1 snk_2000 snk_3700 snk_test0 snk_5000_0 ena_src_200_0 ena_snk_test1 ena_src_400 ena_snk_test0 ena_src_600
*+ avss ena_src_10000_1 dvdd ena_src_10000_0 ena_src_test1 ena_src_test0 ref_sel_vbg ref_in dvss
*.ipin ref_in
*.iopin avss
*.ipin ref_sel_vbg
*.iopin avdd
*.ipin ena_src_test0
*.ipin ena_snk_test0
*.iopin src_test0
*.iopin snk_test0
*.ipin ena_snk_test1
*.iopin snk_test1
*.ipin ena_src_test1
*.iopin src_test1
*.ipin ena_src_10000_0
*.iopin src_10000_0
*.ipin ena_snk_5000_0
*.iopin snk_5000_0
*.ipin ena_src_10000_1
*.iopin src_10000_1
*.ipin ena_snk_5000_1
*.iopin snk_5000_1
*.ipin ena_snk_5000_2
*.iopin snk_5000_2
*.ipin ena_src_600
*.iopin src_600
*.ipin ena_src_400
*.iopin src_400
*.ipin ena_src_200_0
*.iopin src_200_0
*.ipin ena_src_200_1
*.iopin src_200_1
*.ipin ena_src_200_2
*.iopin src_200_2
*.ipin ena_src_100
*.iopin src_100
*.ipin ena_src_50
*.iopin src_50
*.ipin ena_snk_3700
*.iopin snk_3700
*.ipin ena_snk_2000
*.iopin snk_2000
*.ipin vbg
*.ipin ena
*.iopin dvdd
*.iopin dvss
x2[19] net1 ena_3v3 nbias nbias avss bias_nstack
x2[18] net1 ena_3v3 nbias nbias avss bias_nstack
x2[17] net1 ena_3v3 nbias nbias avss bias_nstack
x2[16] net1 ena_3v3 nbias nbias avss bias_nstack
x2[15] net1 ena_3v3 nbias nbias avss bias_nstack
x2[14] net1 ena_3v3 nbias nbias avss bias_nstack
x2[13] net1 ena_3v3 nbias nbias avss bias_nstack
x2[12] net1 ena_3v3 nbias nbias avss bias_nstack
x2[11] net1 ena_3v3 nbias nbias avss bias_nstack
x2[10] net1 ena_3v3 nbias nbias avss bias_nstack
x2[9] net1 ena_3v3 nbias nbias avss bias_nstack
x2[8] net1 ena_3v3 nbias nbias avss bias_nstack
x2[7] net1 ena_3v3 nbias nbias avss bias_nstack
x2[6] net1 ena_3v3 nbias nbias avss bias_nstack
x2[5] net1 ena_3v3 nbias nbias avss bias_nstack
x2[4] net1 ena_3v3 nbias nbias avss bias_nstack
x2[3] net1 ena_3v3 nbias nbias avss bias_nstack
x2[2] net1 ena_3v3 nbias nbias avss bias_nstack
x2[1] net1 ena_3v3 nbias nbias avss bias_nstack
x2[0] net1 ena_3v3 nbias nbias avss bias_nstack
XR3 net1 net15 avss sky130_fd_pr__res_high_po_0p35 L=450 mult=1 m=1
XR4 pcasc ref_in avss sky130_fd_pr__res_high_po_0p35 L=1500 mult=1 m=1
x4 net2 enb_vbg_3v3 net14 nbias avss bias_nstack
x2 avdd pbias pcasc pbias ena_vbg_3v3 avss net2 bias_pstack
x13[1] avdd pbias pcasc net18 enb_test0_3v3 avss src_test0 bias_pstack
x13[0] avdd pbias pcasc net18 enb_test0_3v3 avss src_test0 bias_pstack
x17[1] snk_test0 ena_test0_3v3 net19 nbias avss bias_nstack
x17[0] snk_test0 ena_test0_3v3 net19 nbias avss bias_nstack
x18[1] snk_test1 ena_test1_3v3 net20 nbias avss bias_nstack
x18[0] snk_test1 ena_test1_3v3 net20 nbias avss bias_nstack
x16[1] avdd pbias pcasc net21 enb_test1_3v3 avss src_test1 bias_pstack
x16[0] avdd pbias pcasc net21 enb_test1_3v3 avss src_test1 bias_pstack
x8[199] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[198] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[197] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[196] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[195] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[194] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[193] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[192] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[191] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[190] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[189] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[188] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[187] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[186] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[185] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[184] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[183] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[182] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[181] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[180] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[179] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[178] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[177] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[176] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[175] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[174] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[173] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[172] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[171] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[170] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[169] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[168] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[167] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[166] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[165] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[164] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[163] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[162] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[161] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[160] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[159] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[158] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[157] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[156] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[155] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[154] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[153] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[152] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[151] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[150] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[149] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[148] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[147] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[146] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[145] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[144] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[143] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[142] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[141] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[140] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[139] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[138] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[137] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[136] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[135] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[134] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[133] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[132] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[131] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[130] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[129] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[128] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[127] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[126] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[125] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[124] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[123] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[122] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[121] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[120] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[119] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[118] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[117] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[116] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[115] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[114] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[113] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[112] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[111] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[110] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[109] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[108] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[107] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[106] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[105] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[104] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[103] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[102] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[101] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[100] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[99] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[98] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[97] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[96] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[95] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[94] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[93] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[92] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[91] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[90] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[89] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[88] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[87] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[86] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[85] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[84] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[83] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[82] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[81] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[80] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[79] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[78] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[77] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[76] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[75] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[74] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[73] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[72] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[71] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[70] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[69] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[68] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[67] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[66] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[65] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[64] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[63] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[62] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[61] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[60] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[59] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[58] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[57] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[56] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[55] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[54] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[53] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[52] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[51] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[50] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[49] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[48] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[47] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[46] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[45] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[44] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[43] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[42] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[41] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[40] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[39] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[38] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[37] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[36] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[35] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[34] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[33] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[32] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[31] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[30] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[29] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[28] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[27] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[26] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[25] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[24] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[23] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[22] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[21] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[20] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[19] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[18] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[17] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[16] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[15] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[14] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[13] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[12] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[11] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[10] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[9] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[8] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[7] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[6] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[5] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[4] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[3] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[2] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[1] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x8[0] avdd pbias pcasc net22 enb_10000_0_3v3 avss src_10000_0 bias_pstack
x9[99] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[98] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[97] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[96] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[95] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[94] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[93] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[92] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[91] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[90] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[89] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[88] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[87] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[86] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[85] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[84] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[83] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[82] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[81] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[80] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[79] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[78] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[77] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[76] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[75] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[74] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[73] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[72] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[71] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[70] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[69] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[68] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[67] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[66] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[65] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[64] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[63] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[62] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[61] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[60] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[59] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[58] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[57] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[56] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[55] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[54] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[53] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[52] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[51] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[50] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[49] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[48] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[47] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[46] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[45] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[44] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[43] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[42] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[41] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[40] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[39] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[38] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[37] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[36] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[35] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[34] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[33] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[32] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[31] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[30] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[29] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[28] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[27] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[26] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[25] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[24] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[23] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[22] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[21] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[20] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[19] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[18] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[17] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[16] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[15] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[14] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[13] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[12] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[11] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[10] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[9] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[8] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[7] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[6] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[5] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[4] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[3] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[2] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[1] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x9[0] snk_5000_0 ena_5000_0_3v3 net23 nbias avss bias_nstack
x10[199] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[198] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[197] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[196] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[195] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[194] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[193] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[192] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[191] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[190] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[189] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[188] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[187] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[186] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[185] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[184] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[183] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[182] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[181] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[180] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[179] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[178] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[177] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[176] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[175] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[174] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[173] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[172] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[171] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[170] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[169] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[168] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[167] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[166] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[165] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[164] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[163] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[162] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[161] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[160] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[159] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[158] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[157] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[156] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[155] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[154] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[153] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[152] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[151] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[150] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[149] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[148] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[147] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[146] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[145] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[144] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[143] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[142] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[141] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[140] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[139] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[138] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[137] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[136] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[135] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[134] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[133] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[132] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[131] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[130] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[129] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[128] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[127] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[126] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[125] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[124] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[123] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[122] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[121] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[120] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[119] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[118] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[117] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[116] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[115] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[114] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[113] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[112] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[111] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[110] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[109] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[108] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[107] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[106] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[105] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[104] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[103] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[102] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[101] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[100] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[99] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[98] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[97] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[96] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[95] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[94] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[93] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[92] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[91] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[90] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[89] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[88] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[87] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[86] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[85] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[84] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[83] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[82] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[81] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[80] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[79] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[78] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[77] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[76] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[75] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[74] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[73] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[72] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[71] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[70] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[69] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[68] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[67] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[66] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[65] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[64] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[63] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[62] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[61] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[60] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[59] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[58] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[57] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[56] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[55] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[54] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[53] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[52] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[51] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[50] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[49] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[48] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[47] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[46] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[45] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[44] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[43] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[42] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[41] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[40] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[39] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[38] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[37] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[36] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[35] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[34] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[33] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[32] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[31] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[30] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[29] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[28] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[27] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[26] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[25] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[24] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[23] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[22] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[21] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[20] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[19] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[18] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[17] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[16] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[15] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[14] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[13] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[12] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[11] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[10] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[9] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[8] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[7] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[6] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[5] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[4] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[3] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[2] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[1] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x10[0] avdd pbias pcasc net24 enb_10000_1_3v3 avss src_10000_1 bias_pstack
x1[99] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[98] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[97] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[96] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[95] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[94] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[93] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[92] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[91] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[90] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[89] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[88] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[87] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[86] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[85] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[84] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[83] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[82] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[81] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[80] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[79] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[78] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[77] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[76] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[75] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[74] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[73] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[72] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[71] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[70] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[69] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[68] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[67] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[66] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[65] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[64] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[63] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[62] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[61] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[60] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[59] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[58] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[57] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[56] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[55] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[54] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[53] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[52] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[51] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[50] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[49] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[48] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[47] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[46] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[45] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[44] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[43] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[42] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[41] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[40] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[39] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[38] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[37] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[36] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[35] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[34] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[33] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[32] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[31] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[30] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[29] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[28] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[27] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[26] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[25] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[24] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[23] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[22] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[21] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[20] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[19] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[18] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[17] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[16] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[15] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[14] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[13] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[12] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[11] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[10] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[9] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[8] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[7] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[6] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[5] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[4] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[3] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[2] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[1] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x1[0] snk_5000_1 ena_5000_1_3v3 net25 nbias avss bias_nstack
x3[99] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[98] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[97] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[96] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[95] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[94] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[93] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[92] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[91] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[90] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[89] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[88] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[87] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[86] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[85] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[84] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[83] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[82] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[81] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[80] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[79] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[78] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[77] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[76] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[75] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[74] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[73] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[72] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[71] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[70] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[69] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[68] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[67] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[66] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[65] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[64] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[63] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[62] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[61] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[60] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[59] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[58] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[57] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[56] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[55] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[54] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[53] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[52] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[51] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[50] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[49] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[48] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[47] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[46] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[45] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[44] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[43] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[42] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[41] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[40] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[39] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[38] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[37] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[36] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[35] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[34] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[33] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[32] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[31] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[30] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[29] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[28] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[27] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[26] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[25] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[24] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[23] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[22] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[21] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[20] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[19] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[18] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[17] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[16] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[15] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[14] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[13] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[12] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[11] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[10] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[9] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[8] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[7] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[6] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[5] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[4] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[3] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[2] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[1] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x3[0] snk_5000_2 ena_5000_2_3v3 net26 nbias avss bias_nstack
x4[11] avdd pbias pcasc net27 enb_600_3v3 avss src_600 bias_pstack
x4[10] avdd pbias pcasc net27 enb_600_3v3 avss src_600 bias_pstack
x4[9] avdd pbias pcasc net27 enb_600_3v3 avss src_600 bias_pstack
x4[8] avdd pbias pcasc net27 enb_600_3v3 avss src_600 bias_pstack
x4[7] avdd pbias pcasc net27 enb_600_3v3 avss src_600 bias_pstack
x4[6] avdd pbias pcasc net27 enb_600_3v3 avss src_600 bias_pstack
x4[5] avdd pbias pcasc net27 enb_600_3v3 avss src_600 bias_pstack
x4[4] avdd pbias pcasc net27 enb_600_3v3 avss src_600 bias_pstack
x4[3] avdd pbias pcasc net27 enb_600_3v3 avss src_600 bias_pstack
x4[2] avdd pbias pcasc net27 enb_600_3v3 avss src_600 bias_pstack
x4[1] avdd pbias pcasc net27 enb_600_3v3 avss src_600 bias_pstack
x4[0] avdd pbias pcasc net27 enb_600_3v3 avss src_600 bias_pstack
x5[7] avdd pbias pcasc net28 enb_400_3v3 avss src_400 bias_pstack
x5[6] avdd pbias pcasc net28 enb_400_3v3 avss src_400 bias_pstack
x5[5] avdd pbias pcasc net28 enb_400_3v3 avss src_400 bias_pstack
x5[4] avdd pbias pcasc net28 enb_400_3v3 avss src_400 bias_pstack
x5[3] avdd pbias pcasc net28 enb_400_3v3 avss src_400 bias_pstack
x5[2] avdd pbias pcasc net28 enb_400_3v3 avss src_400 bias_pstack
x5[1] avdd pbias pcasc net28 enb_400_3v3 avss src_400 bias_pstack
x5[0] avdd pbias pcasc net28 enb_400_3v3 avss src_400 bias_pstack
x6[3] avdd pbias pcasc net29 enb_200_0_3v3 avss src_200_0 bias_pstack
x6[2] avdd pbias pcasc net29 enb_200_0_3v3 avss src_200_0 bias_pstack
x6[1] avdd pbias pcasc net29 enb_200_0_3v3 avss src_200_0 bias_pstack
x6[0] avdd pbias pcasc net29 enb_200_0_3v3 avss src_200_0 bias_pstack
x7[3] avdd pbias pcasc net30 enb_200_1_3v3 avss src_200_1 bias_pstack
x7[2] avdd pbias pcasc net30 enb_200_1_3v3 avss src_200_1 bias_pstack
x7[1] avdd pbias pcasc net30 enb_200_1_3v3 avss src_200_1 bias_pstack
x7[0] avdd pbias pcasc net30 enb_200_1_3v3 avss src_200_1 bias_pstack
x11[3] avdd pbias pcasc net31 enb_200_2_3v3 avss src_200_2 bias_pstack
x11[2] avdd pbias pcasc net31 enb_200_2_3v3 avss src_200_2 bias_pstack
x11[1] avdd pbias pcasc net31 enb_200_2_3v3 avss src_200_2 bias_pstack
x11[0] avdd pbias pcasc net31 enb_200_2_3v3 avss src_200_2 bias_pstack
x12[1] avdd pbias pcasc net32 enb_100_3v3 avss src_100 bias_pstack
x12[0] avdd pbias pcasc net32 enb_100_3v3 avss src_100 bias_pstack
x13 avdd pbias pcasc net33 enb_50_3v3 avss src_50 bias_pstack
x14[74] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[73] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[72] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[71] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[70] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[69] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[68] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[67] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[66] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[65] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[64] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[63] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[62] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[61] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[60] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[59] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[58] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[57] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[56] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[55] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[54] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[53] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[52] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[51] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[50] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[49] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[48] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[47] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[46] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[45] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[44] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[43] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[42] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[41] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[40] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[39] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[38] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[37] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[36] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[35] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[34] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[33] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[32] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[31] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[30] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[29] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[28] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[27] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[26] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[25] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[24] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[23] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[22] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[21] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[20] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[19] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[18] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[17] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[16] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[15] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[14] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[13] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[12] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[11] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[10] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[9] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[8] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[7] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[6] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[5] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[4] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[3] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[2] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[1] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x14[0] snk_3700 ena_3700_3v3 net34 nbias avss bias_nstack
x15[39] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[38] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[37] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[36] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[35] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[34] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[33] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[32] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[31] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[30] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[29] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[28] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[27] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[26] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[25] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[24] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[23] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[22] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[21] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[20] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[19] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[18] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[17] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[16] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[15] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[14] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[13] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[12] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[11] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[10] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[9] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[8] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[7] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[6] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[5] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[4] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[3] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[2] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[1] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x15[0] snk_2000 enb_2000_3v3 net35 nbias avss bias_nstack
x1 ref_sel_vbg dvdd dvss dvss avdd avdd ena_vbg_3v3 sky130_fd_sc_hvl__lsbuflv2hv_1
x5 ena_snk_2000 dvdd dvss dvss avdd avdd enb_2000_3v3 sky130_fd_sc_hvl__lsbuflv2hv_1
x6 ena_snk_3700 dvdd dvss dvss avdd avdd ena_3700_3v3 sky130_fd_sc_hvl__lsbuflv2hv_1
x7 ena_snk_5000_2 dvdd dvss dvss avdd avdd ena_5000_2_3v3 sky130_fd_sc_hvl__lsbuflv2hv_1
x8 ena_snk_5000_1 dvdd dvss dvss avdd avdd ena_5000_1_3v3 sky130_fd_sc_hvl__lsbuflv2hv_1
x9 ena_snk_5000_0 dvdd dvss dvss avdd avdd ena_5000_0_3v3 sky130_fd_sc_hvl__lsbuflv2hv_1
x10 ena_snk_test1 dvdd dvss dvss avdd avdd ena_test1_3v3 sky130_fd_sc_hvl__lsbuflv2hv_1
x11 ena_snk_test0 dvdd dvss dvss avdd avdd ena_test0_3v3 sky130_fd_sc_hvl__lsbuflv2hv_1
x12 ena_src_50 dvdd dvss dvss avdd avdd net13 sky130_fd_sc_hvl__lsbuflv2hv_1
x14 ena_src_100 dvdd dvss dvss avdd avdd net12 sky130_fd_sc_hvl__lsbuflv2hv_1
x15 ena_src_200_2 dvdd dvss dvss avdd avdd net11 sky130_fd_sc_hvl__lsbuflv2hv_1
x16 ena_src_200_1 dvdd dvss dvss avdd avdd net10 sky130_fd_sc_hvl__lsbuflv2hv_1
x17 ena_src_200_0 dvdd dvss dvss avdd avdd net9 sky130_fd_sc_hvl__lsbuflv2hv_1
x18 ena_src_400 dvdd dvss dvss avdd avdd net8 sky130_fd_sc_hvl__lsbuflv2hv_1
x19 ena_src_600 dvdd dvss dvss avdd avdd net7 sky130_fd_sc_hvl__lsbuflv2hv_1
x20 ena_src_10000_1 dvdd dvss dvss avdd avdd net6 sky130_fd_sc_hvl__lsbuflv2hv_1
x21 ena_src_10000_0 dvdd dvss dvss avdd avdd net5 sky130_fd_sc_hvl__lsbuflv2hv_1
x22 ena_src_test1 dvdd dvss dvss avdd avdd net4 sky130_fd_sc_hvl__lsbuflv2hv_1
x23 ena_src_test0 dvdd dvss dvss avdd avdd net3 sky130_fd_sc_hvl__lsbuflv2hv_1
x24 ena_vbg_3v3 dvss dvss avdd avdd enb_vbg_3v3 sky130_fd_sc_hvl__inv_2
x25 net13 dvss dvss avdd avdd enb_50_3v3 sky130_fd_sc_hvl__inv_2
x26 net12 dvss dvss avdd avdd enb_100_3v3 sky130_fd_sc_hvl__inv_2
x27 net11 dvss dvss avdd avdd enb_200_2_3v3 sky130_fd_sc_hvl__inv_2
x28 net10 dvss dvss avdd avdd enb_200_1_3v3 sky130_fd_sc_hvl__inv_2
x29 net9 dvss dvss avdd avdd enb_200_0_3v3 sky130_fd_sc_hvl__inv_2
x30 net8 dvss dvss avdd avdd enb_400_3v3 sky130_fd_sc_hvl__inv_2
x31 net7 dvss dvss avdd avdd enb_600_3v3 sky130_fd_sc_hvl__inv_2
x32 net6 dvss dvss avdd avdd enb_10000_1_3v3 sky130_fd_sc_hvl__inv_2
x33 net5 dvss dvss avdd avdd enb_10000_0_3v3 sky130_fd_sc_hvl__inv_2
x34 net4 dvss dvss avdd avdd enb_test1_3v3 sky130_fd_sc_hvl__inv_2
x35 net3 dvss dvss avdd avdd enb_test0_3v3 sky130_fd_sc_hvl__inv_2
x3 avdd pbias vbg vfb nbias avss ena_vbg_3v3 bias_amp
XR1 avss net17 avss sky130_fd_pr__res_high_po_0p35 L=1328 mult=1 m=1
XC1 pbias vfb sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=8 m=8
x36 ena dvdd dvss dvss avdd avdd ena_3v3 sky130_fd_sc_hvl__lsbuflv2hv_1
x37 ena_3v3 dvss dvss avdd avdd enb_3v3 sky130_fd_sc_hvl__inv_2
* noconn #net14
* noconn #net19
* noconn #net18
* noconn #net21
* noconn #net20
* noconn #net23
* noconn #net22
* noconn #net25
* noconn #net24
* noconn #net27
* noconn #net26
* noconn #net34
* noconn #net28
* noconn #net35
* noconn #net29
* noconn #net30
* noconn #net31
* noconn #net32
* noconn #net33
XR2 net15 pcasc avss sky130_fd_pr__res_high_po_0p35 L=450 mult=1 m=1
Vmeas net16 net17 0
.save i(vmeas)
x19[11] avdd pbias pcasc vfb enb_vbg_3v3 avss net16 bias_pstack
x19[10] avdd pbias pcasc vfb enb_vbg_3v3 avss net16 bias_pstack
x19[9] avdd pbias pcasc vfb enb_vbg_3v3 avss net16 bias_pstack
x19[8] avdd pbias pcasc vfb enb_vbg_3v3 avss net16 bias_pstack
x19[7] avdd pbias pcasc vfb enb_vbg_3v3 avss net16 bias_pstack
x19[6] avdd pbias pcasc vfb enb_vbg_3v3 avss net16 bias_pstack
x19[5] avdd pbias pcasc vfb enb_vbg_3v3 avss net16 bias_pstack
x19[4] avdd pbias pcasc vfb enb_vbg_3v3 avss net16 bias_pstack
x19[3] avdd pbias pcasc vfb enb_vbg_3v3 avss net16 bias_pstack
x19[2] avdd pbias pcasc vfb enb_vbg_3v3 avss net16 bias_pstack
x19[1] avdd pbias pcasc vfb enb_vbg_3v3 avss net16 bias_pstack
x19[0] avdd pbias pcasc vfb enb_vbg_3v3 avss net16 bias_pstack
**.ends

* expanding   symbol:  bias_nstack.sym # of pins=5
** sym_path: /home/tim/gits/sky130_ef_ip__biasgen/xschem/bias_nstack.sym
** sch_path: /home/tim/gits/sky130_ef_ip__biasgen/xschem/bias_nstack.sch
.subckt bias_nstack itail ena vcasc nbias avss
*.iopin avss
*.ipin ena
*.ipin nbias
*.iopin itail
*.iopin vcasc
XM3 net1 nbias avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 vcasc nbias net1 avss sky130_fd_pr__nfet_05v0_nvt L=1 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 itail ena vcasc avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XD1 avss ena sky130_fd_pr__diode_pw2nd_05v5 area=2.025e11 perim=1.8e6
.ends


* expanding   symbol:  bias_pstack.sym # of pins=7
** sym_path: /home/tim/gits/sky130_ef_ip__biasgen/xschem/bias_pstack.sym
** sch_path: /home/tim/gits/sky130_ef_ip__biasgen/xschem/bias_pstack.sch
.subckt bias_pstack avdd pbias pcasc vcasc enb avss itail
*.iopin avdd
*.iopin itail
*.ipin enb
*.ipin pcasc
*.iopin vcasc
*.ipin pbias
*.iopin avss
XM13 net1 pbias avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM18 itail enb vcasc avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM14 vcasc pcasc net1 avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XD1 avss enb sky130_fd_pr__diode_pw2nd_05v5 area=2.025e11 perim=1.8e6
.ends


* expanding   symbol:  bias_amp.sym # of pins=7
** sym_path: /home/tim/gits/sky130_ef_ip__biasgen/xschem/bias_amp.sym
** sch_path: /home/tim/gits/sky130_ef_ip__biasgen/xschem/bias_amp.sch
.subckt bias_amp avdd out inn inp nbias avss ena
*.ipin inp
*.ipin nbias
*.ipin inn
*.opin out
*.iopin avdd
*.iopin avss
*.ipin ena
XM1 net2 nbias avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 out net1 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 net1 net1 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net1 inp vcom avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=4 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 out inn vcom avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=4 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 vcom ena net2 avss sky130_fd_pr__nfet_05v0_nvt L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
