magic
tech sky130A
magscale 1 2
timestamp 1715390562
<< dnwell >>
rect -896 -5634 248954 2218
<< nwell >>
rect -1005 2012 249063 2327
rect -1005 -5428 -690 2012
rect 248748 -5428 249063 2012
rect -1005 -5743 249063 -5428
<< pwell >>
rect -453 -5169 -383 -4737
rect 15100 -5428 15188 -5406
<< mvpsubdiff >>
rect -1125 2417 -1065 2451
rect 249123 2417 249183 2451
rect -1125 2391 -1091 2417
rect 249149 2391 249183 2417
rect -1125 -5855 -1091 -5829
rect 249149 -5855 249183 -5829
rect -1125 -5889 -1065 -5855
rect 249123 -5889 249183 -5855
<< mvnsubdiff >>
rect -939 2241 248997 2261
rect -939 2207 -859 2241
rect 248917 2207 248997 2241
rect -939 2187 248997 2207
rect -939 2181 -865 2187
rect -939 -5597 -919 2181
rect -885 -5597 -865 2181
rect -939 -5603 -865 -5597
rect 248923 2181 248997 2187
rect 248923 -5597 248943 2181
rect 248977 -5597 248997 2181
rect 248923 -5603 248997 -5597
rect -939 -5623 248997 -5603
rect -939 -5657 -859 -5623
rect 248917 -5657 248997 -5623
rect -939 -5677 248997 -5657
<< mvpsubdiffcont >>
rect -1065 2417 249123 2451
rect -1125 -5829 -1091 2391
rect 249149 -5829 249183 2391
rect -1065 -5889 249123 -5855
<< mvnsubdiffcont >>
rect -859 2207 248917 2241
rect -919 -5597 -885 2181
rect 248943 -5597 248977 2181
rect -859 -5657 248917 -5623
<< locali >>
rect -1125 2417 -1065 2451
rect 249123 2417 249183 2451
rect -1125 2402 249183 2417
rect -1125 2391 249085 2402
rect -1091 2318 249085 2391
rect -1091 -3629 -1023 2318
rect -1050 -5711 -1023 -3629
rect -919 2207 -859 2241
rect 248917 2207 248977 2241
rect -919 2181 248977 2207
rect -885 2176 248943 2181
rect -885 2022 248853 2176
rect -885 -5444 -751 2022
rect 248806 -5444 248853 2022
rect -885 -5597 248853 -5444
rect -919 -5601 248853 -5597
rect 248912 -5597 248943 2176
rect 248912 -5601 248977 -5597
rect -919 -5623 248977 -5601
rect -919 -5657 -859 -5623
rect 248917 -5657 248977 -5623
rect -1091 -5743 -1023 -5711
rect 249041 -5743 249085 2318
rect -1091 -5829 249085 -5743
rect -1125 -5830 249085 -5829
rect -1125 -5874 -1098 -5830
rect 249032 -5839 249085 -5830
rect 249137 2391 249183 2402
rect 249137 -5829 249149 2391
rect 249137 -5839 249183 -5829
rect 249032 -5855 249183 -5839
rect -1125 -5889 -1065 -5874
rect 249123 -5889 249183 -5855
<< viali >>
rect -1099 -5711 -1091 -3629
rect -1091 -5711 -1050 -3629
rect 248853 -5601 248912 2176
rect -1098 -5855 249032 -5830
rect 249085 -5839 249137 2402
rect -1098 -5874 -1065 -5855
rect -1065 -5874 249032 -5855
<< metal1 >>
rect 249057 2402 249173 2444
rect 248818 2176 248956 2227
rect -583 1818 12861 1829
rect -583 1766 -550 1818
rect 12825 1766 12861 1818
rect -583 1754 12861 1766
rect -583 1431 -383 1663
rect -902 1231 -383 1431
rect -287 1231 -51 1663
rect 45 1231 281 1663
rect 377 1231 613 1663
rect 709 1231 945 1663
rect 1041 1231 1277 1663
rect 1373 1231 1609 1663
rect 1705 1231 1941 1663
rect 2037 1231 2273 1663
rect 2369 1231 2605 1663
rect 2701 1231 2937 1663
rect 3033 1231 3269 1663
rect 3365 1231 3601 1663
rect 3697 1231 3933 1663
rect 4029 1231 4265 1663
rect 4361 1231 4597 1663
rect 4693 1231 4929 1663
rect 5025 1231 5261 1663
rect 5357 1231 5593 1663
rect 5689 1231 5925 1663
rect 6021 1231 6257 1663
rect 6353 1231 6589 1663
rect 6685 1231 6921 1663
rect 7017 1231 7253 1663
rect 7349 1231 7585 1663
rect -1125 -3629 -1023 -3590
rect -1125 -3754 -1099 -3629
rect -1127 -5313 -1099 -3754
rect -1125 -5711 -1099 -5313
rect -1050 -3754 -1023 -3629
rect -1050 -3774 -681 -3754
rect -1050 -5294 -860 -3774
rect -704 -5294 -681 -3774
rect -1050 -5313 -681 -5294
rect -589 -4869 -537 1069
rect 7681 577 7917 1663
rect 8013 1231 8249 1663
rect 8345 1231 8581 1663
rect 8677 1231 8913 1663
rect 9009 1231 9245 1663
rect 9341 1231 9577 1663
rect 9673 1231 9909 1663
rect 10005 1231 10241 1663
rect 10337 1231 10573 1663
rect 10669 1231 10905 1663
rect 11001 1231 11237 1663
rect 11333 1231 11569 1663
rect 11665 1231 11901 1663
rect 11997 1231 12233 1663
rect 12329 1231 12565 1663
rect 12660 1371 12861 1663
rect 12660 1231 13108 1371
rect 7681 328 7917 343
rect 12821 -1873 12873 -1859
rect 12821 -2125 12873 -2111
rect 12968 -3739 13108 1231
rect 248818 -54 248853 2176
rect 248912 -54 248956 2176
rect 46785 -427 46853 -318
rect 46635 -661 46785 -459
rect 46635 -705 46853 -661
rect 248818 -1696 248833 -54
rect 248940 -1696 248956 -54
rect 36120 -2897 36182 -2882
rect 36120 -3228 36182 -3135
rect 36654 -2897 36716 -2882
rect 36654 -3228 36716 -3135
rect 37188 -2897 37250 -2882
rect 37188 -3228 37250 -3135
rect 37722 -2897 37784 -2882
rect 37722 -3228 37784 -3135
rect 38256 -2897 38318 -2882
rect 38256 -3228 38318 -3135
rect 38790 -2897 38852 -2882
rect 38790 -3228 38852 -3135
rect 39324 -2897 39386 -2882
rect 39324 -3228 39386 -3135
rect 39858 -2897 39920 -2882
rect 39858 -3228 39920 -3135
rect 40392 -2897 40454 -2882
rect 40392 -3228 40454 -3135
rect 40926 -2897 40988 -2882
rect 40926 -3228 40988 -3135
rect 41460 -2897 41522 -2882
rect 41460 -3228 41522 -3135
rect 41994 -2897 42056 -2882
rect 41994 -3228 42056 -3135
rect 42528 -2897 42590 -2882
rect 42528 -3228 42590 -3135
rect 43062 -2897 43124 -2882
rect 43062 -3228 43124 -3135
rect 43596 -2897 43658 -2882
rect 43596 -3228 43658 -3135
rect 44130 -2897 44192 -2882
rect 44130 -3228 44192 -3135
rect 44664 -2897 44726 -2882
rect 44664 -3228 44726 -3135
rect 45198 -2897 45260 -2882
rect 45198 -3228 45260 -3135
rect 45732 -2897 45794 -2882
rect 45732 -3228 45794 -3135
rect 46266 -2897 46328 -2882
rect 46266 -3228 46328 -3135
rect 36320 -3881 36384 -3871
rect 36320 -4194 36384 -4119
rect 36854 -3881 36918 -3871
rect 36854 -4194 36918 -4119
rect 37388 -3881 37452 -3871
rect 37388 -4194 37452 -4119
rect 37922 -3881 37986 -3871
rect 37922 -4194 37986 -4119
rect 38456 -3881 38520 -3871
rect 38456 -4194 38520 -4119
rect 38990 -3881 39054 -3871
rect 38990 -4194 39054 -4119
rect 39516 -3881 39588 -3871
rect 39516 -4194 39588 -4119
rect 40050 -3881 40122 -3871
rect 40050 -4194 40122 -4119
rect 40584 -3881 40656 -3871
rect 40584 -4194 40656 -4119
rect 41118 -3881 41190 -3871
rect 41118 -4194 41190 -4119
rect 41652 -3881 41724 -3871
rect 41652 -4194 41724 -4119
rect 42186 -3881 42258 -3871
rect 42186 -4194 42258 -4119
rect 42720 -3881 42792 -3871
rect 42720 -4194 42792 -4119
rect 43254 -3881 43326 -3871
rect 43254 -4194 43326 -4119
rect 43788 -3881 43852 -3871
rect 43788 -4194 43852 -4119
rect 44322 -3881 44386 -3871
rect 44322 -4194 44386 -4119
rect 44856 -3881 44920 -3871
rect 44856 -4194 44920 -4119
rect 45390 -3881 45454 -3871
rect 45390 -4194 45454 -4119
rect 45924 -3881 45988 -3871
rect 45924 -4194 45988 -4119
rect 12968 -4262 13108 -4225
rect -589 -5305 -537 -5107
rect -453 -5169 -217 -4737
rect -121 -5169 115 -4737
rect 211 -5169 447 -4737
rect 543 -5169 779 -4737
rect 875 -5169 1111 -4737
rect 1207 -5169 1443 -4737
rect 1539 -5169 1775 -4737
rect 1871 -5169 2107 -4737
rect 2203 -5169 2439 -4737
rect 2535 -5169 2771 -4737
rect 2867 -5169 3103 -4737
rect 3199 -5169 3435 -4737
rect 3531 -5169 3767 -4737
rect 3863 -5169 4099 -4737
rect 4195 -5169 4431 -4737
rect 4527 -5169 4763 -4737
rect 4859 -5169 5095 -4737
rect 5191 -5169 5427 -4737
rect 5523 -5169 5759 -4737
rect 5855 -5169 6091 -4737
rect 6187 -5169 6423 -4737
rect 6519 -5169 6755 -4737
rect 6851 -5169 7087 -4737
rect 7183 -5169 7419 -4737
rect 7515 -5169 7751 -4737
rect 7847 -5169 8083 -4737
rect 8179 -5169 8415 -4737
rect 8511 -5169 8747 -4737
rect 8843 -5169 9079 -4737
rect 9175 -5169 9411 -4737
rect 9507 -5169 9743 -4737
rect 9839 -5169 10075 -4737
rect 10171 -5169 10407 -4737
rect 10503 -5169 10739 -4737
rect 10835 -5169 11071 -4737
rect 11167 -5169 11403 -4737
rect 11499 -5169 11735 -4737
rect 11831 -5169 12067 -4737
rect 12163 -5169 12399 -4737
rect 12495 -5169 12731 -4737
rect 12821 -5305 12867 -4575
rect -1050 -5711 -1023 -5313
rect 36494 -5532 36548 -5504
rect 37028 -5532 37082 -5504
rect 37562 -5532 37616 -5504
rect 38096 -5532 38150 -5504
rect 38630 -5532 38684 -5504
rect 39164 -5532 39218 -5504
rect 39698 -5532 39752 -5504
rect 40232 -5532 40286 -5504
rect 40766 -5532 40820 -5504
rect 41300 -5532 41354 -5504
rect 41834 -5532 41888 -5504
rect 42368 -5532 42422 -5504
rect 42902 -5532 42956 -5504
rect 43436 -5532 43490 -5504
rect 43970 -5532 44024 -5504
rect 44504 -5532 44558 -5504
rect 45038 -5532 45092 -5504
rect 45572 -5532 45626 -5504
rect 46106 -5532 46160 -5504
rect 46640 -5532 46694 -5504
rect 248818 -5601 248853 -1696
rect 248912 -5601 248956 -1696
rect 248818 -5648 248956 -5601
rect -1125 -5811 -1023 -5711
rect 249057 -5811 249085 2402
rect -1125 -5830 249085 -5811
rect -1125 -5874 -1098 -5830
rect 249032 -5839 249085 -5830
rect 249137 -5839 249173 2402
rect 249032 -5874 249173 -5839
rect -1125 -5889 249173 -5874
<< via1 >>
rect 46639 2384 46693 2616
rect -550 1766 12825 1818
rect -860 -5294 -704 -3774
rect 7681 343 7917 577
rect 12821 -2111 12873 -1873
rect 46480 677 46549 1236
rect 46785 -661 46853 -427
rect 248833 -1696 248853 -54
rect 248853 -1696 248912 -54
rect 248912 -1696 248940 -54
rect 36120 -3135 36182 -2897
rect 36654 -3135 36716 -2897
rect 37188 -3135 37250 -2897
rect 37722 -3135 37784 -2897
rect 38256 -3135 38318 -2897
rect 38790 -3135 38852 -2897
rect 39324 -3135 39386 -2897
rect 39858 -3135 39920 -2897
rect 40392 -3135 40454 -2897
rect 40926 -3135 40988 -2897
rect 41460 -3135 41522 -2897
rect 41994 -3135 42056 -2897
rect 42528 -3135 42590 -2897
rect 43062 -3135 43124 -2897
rect 43596 -3135 43658 -2897
rect 44130 -3135 44192 -2897
rect 44664 -3135 44726 -2897
rect 45198 -3135 45260 -2897
rect 45732 -3135 45794 -2897
rect 46266 -3135 46328 -2897
rect 12968 -4225 13108 -3739
rect 36320 -4119 36384 -3881
rect 36854 -4119 36918 -3881
rect 37388 -4119 37452 -3881
rect 37922 -4119 37986 -3881
rect 38456 -4119 38520 -3881
rect 38990 -4119 39054 -3881
rect 39516 -4119 39588 -3881
rect 40050 -4119 40122 -3881
rect 40584 -4119 40656 -3881
rect 41118 -4119 41190 -3881
rect 41652 -4119 41724 -3881
rect 42186 -4119 42258 -3881
rect 42720 -4119 42792 -3881
rect 43254 -4119 43326 -3881
rect 43788 -4119 43852 -3881
rect 44322 -4119 44386 -3881
rect 44856 -4119 44920 -3881
rect 45390 -4119 45454 -3881
rect 45924 -4119 45988 -3881
rect -589 -5107 -537 -4869
rect 46474 -4774 46562 -4207
rect 36494 -5504 36548 -5316
rect 37028 -5504 37082 -5316
rect 37562 -5504 37616 -5316
rect 38096 -5504 38150 -5316
rect 38630 -5504 38684 -5316
rect 39164 -5504 39218 -5316
rect 39698 -5504 39752 -5316
rect 40232 -5504 40286 -5316
rect 40766 -5504 40820 -5316
rect 41300 -5504 41354 -5316
rect 41834 -5504 41888 -5316
rect 42368 -5504 42422 -5316
rect 42902 -5504 42956 -5316
rect 43436 -5504 43490 -5316
rect 43970 -5504 44024 -5316
rect 44504 -5504 44558 -5316
rect 45038 -5504 45092 -5316
rect 45572 -5504 45626 -5316
rect 46106 -5504 46160 -5316
rect 46640 -5504 46694 -5316
<< metal2 >>
rect 46562 2616 46730 2884
rect 13336 2382 13479 2614
rect 13685 2382 13944 2614
rect 14389 2382 46295 2614
rect 46381 2382 46390 2614
rect 46562 2384 46639 2616
rect 46693 2384 46730 2616
rect 13522 2075 13815 2307
rect 14021 2075 14120 2307
rect 14389 2075 46297 2307
rect 46383 2075 46394 2307
rect 46562 2065 46730 2384
rect 46767 2382 46777 2614
rect 46863 2382 54573 2614
rect 54892 2382 121309 2614
rect 121711 2382 164959 2614
rect 165286 2382 228205 2614
rect 228479 2382 232127 2614
rect 232454 2382 234545 2614
rect 234895 2382 237387 2614
rect 237714 2382 238975 2614
rect 239264 2382 240557 2614
rect 240884 2382 241222 2614
rect 241410 2382 242649 2614
rect 242976 2382 243315 2614
rect 243550 2382 244741 2614
rect 245068 2382 245522 2614
rect 245654 2382 246293 2614
rect 246620 2382 246634 2614
rect 246706 2382 246722 2614
rect 246894 2382 246928 2614
rect 247231 2382 247403 2614
rect 247620 2382 247838 2614
rect 46766 2075 46777 2307
rect 46863 2075 53688 2307
rect 53871 2075 121510 2307
rect 121890 2075 164064 2307
rect 164249 2075 228352 2307
rect 228651 2075 231232 2307
rect 231417 2075 234693 2307
rect 234922 2075 236492 2307
rect 236677 2075 239053 2307
rect 239342 2075 239662 2307
rect 239847 2075 241314 2307
rect 241446 2075 241754 2307
rect 241939 2075 243315 2307
rect 243550 2075 243846 2307
rect 244031 2075 245522 2307
rect 245654 2075 245938 2307
rect 246123 2075 246583 2307
rect 246706 2075 247064 2307
rect 247249 2075 247274 2307
rect 247418 2075 247747 2307
rect 247922 2075 248017 2307
rect -900 1818 12943 1912
rect -900 1766 -550 1818
rect 12825 1766 12943 1818
rect -900 1674 12943 1766
rect 13184 1674 248341 1912
rect -671 1343 13193 1577
rect 248333 1343 248380 1577
rect 248635 1343 248664 1577
rect 46480 1236 46549 1245
rect 46480 668 46549 677
rect -656 343 7681 577
rect 7917 343 248341 577
rect 12960 342 13191 343
rect 248804 -54 248973 -32
rect 13187 -661 46785 -427
rect 46853 -661 248341 -427
rect 248333 -1715 248379 -1481
rect 248634 -1715 248663 -1481
rect 248804 -1696 248833 -54
rect 248940 -1696 248973 -54
rect 248804 -1715 248973 -1696
rect 12811 -2111 12821 -1873
rect 12873 -2111 12944 -1873
rect 13185 -1892 14284 -1873
rect 13185 -1976 13323 -1892
rect 13185 -2111 14284 -1976
rect 13228 -3135 36120 -2897
rect 36182 -3135 36654 -2897
rect 36716 -3135 37188 -2897
rect 37250 -3135 37722 -2897
rect 37784 -3135 38256 -2897
rect 38318 -3135 38790 -2897
rect 38852 -3135 39324 -2897
rect 39386 -3135 39858 -2897
rect 39920 -3135 40392 -2897
rect 40454 -3135 40926 -2897
rect 40988 -3135 41460 -2897
rect 41522 -3135 41994 -2897
rect 42056 -3135 42528 -2897
rect 42590 -3135 43062 -2897
rect 43124 -3135 43596 -2897
rect 43658 -3135 44130 -2897
rect 44192 -3135 44664 -2897
rect 44726 -3135 45198 -2897
rect 45260 -3135 45732 -2897
rect 45794 -3135 46266 -2897
rect 46328 -3135 248322 -2897
rect -1127 -3774 -681 -3754
rect -1127 -5294 -860 -3774
rect -704 -5294 -681 -3774
rect 12956 -4225 12968 -3739
rect 13108 -3881 13119 -3739
rect 13108 -4119 36320 -3881
rect 36384 -4119 36854 -3881
rect 36918 -4119 37388 -3881
rect 37452 -4119 37922 -3881
rect 37986 -4119 38456 -3881
rect 38520 -4119 38990 -3881
rect 39054 -4119 39516 -3881
rect 39588 -4119 40050 -3881
rect 40122 -4119 40584 -3881
rect 40656 -4119 41118 -3881
rect 41190 -4119 41652 -3881
rect 41724 -4119 42186 -3881
rect 42258 -4119 42720 -3881
rect 42792 -4119 43254 -3881
rect 43326 -4119 43788 -3881
rect 43852 -4119 44322 -3881
rect 44386 -4119 44856 -3881
rect 44920 -4119 45390 -3881
rect 45454 -4119 45924 -3881
rect 45988 -4119 248314 -3881
rect 13108 -4225 13119 -4119
rect 12956 -4226 13119 -4225
rect 46474 -4207 46562 -4198
rect 46474 -4783 46562 -4774
rect -612 -5107 -589 -4869
rect -537 -5107 12944 -4869
rect 13185 -5107 248322 -4869
rect -1127 -5313 -681 -5294
rect 12915 -5504 12944 -5316
rect 13070 -5504 14125 -5316
rect 14193 -5504 23221 -5316
rect 23406 -5504 35508 -5316
rect 35572 -5504 36494 -5316
rect 36548 -5504 37028 -5316
rect 37082 -5504 37562 -5316
rect 37616 -5504 38096 -5316
rect 38150 -5504 38630 -5316
rect 38684 -5504 39164 -5316
rect 39218 -5504 39698 -5316
rect 39752 -5504 40232 -5316
rect 40286 -5504 40766 -5316
rect 40820 -5504 41300 -5316
rect 41354 -5504 41834 -5316
rect 41888 -5504 42368 -5316
rect 42422 -5504 42902 -5316
rect 42956 -5504 43436 -5316
rect 43490 -5504 43970 -5316
rect 44024 -5504 44504 -5316
rect 44558 -5504 45038 -5316
rect 45092 -5504 45572 -5316
rect 45626 -5504 46106 -5316
rect 46160 -5504 46640 -5316
rect 46694 -5504 46860 -5316
rect 47157 -5504 69528 -5316
rect 69713 -5504 100124 -5316
rect 100508 -5504 122021 -5316
rect 122206 -5504 153530 -5316
rect 153913 -5504 174621 -5316
rect 174806 -5504 206913 -5316
rect 207335 -5504 230729 -5316
rect 230914 -5504 246964 -5316
rect 247415 -5504 247793 -5316
rect 247910 -5504 248025 -5316
rect 13355 -5760 13541 -5572
rect 13741 -5760 13965 -5572
rect 14412 -5760 24116 -5572
rect 24443 -5760 35340 -5572
rect 35572 -5590 35672 -5504
rect 35472 -5790 35672 -5590
rect 35758 -5760 46004 -5572
rect 46436 -5760 46528 -5572
rect 46986 -5760 70423 -5572
rect 70750 -5760 99970 -5572
rect 100354 -5760 122916 -5572
rect 123243 -5760 153382 -5572
rect 153765 -5760 175516 -5572
rect 175843 -5760 206747 -5572
rect 207169 -5760 231624 -5572
rect 231951 -5760 246806 -5572
rect 247250 -5760 247405 -5572
rect 247587 -5760 247860 -5572
<< via2 >>
rect 13479 2382 13685 2614
rect 46295 2382 46381 2614
rect 13815 2075 14021 2307
rect 46297 2075 46383 2307
rect 46777 2382 46863 2614
rect 54573 2382 54892 2614
rect 164959 2382 165286 2614
rect 232127 2382 232454 2614
rect 237387 2382 237714 2614
rect 240557 2382 240884 2614
rect 242649 2382 242976 2614
rect 244741 2382 245068 2614
rect 246293 2382 246620 2614
rect 246722 2382 246894 2614
rect 247403 2382 247620 2614
rect 46777 2075 46863 2307
rect 53688 2075 53871 2307
rect 164064 2075 164249 2307
rect 231232 2075 231417 2307
rect 236492 2075 236677 2307
rect 239662 2075 239847 2307
rect 241754 2075 241939 2307
rect 243846 2075 244031 2307
rect 245938 2075 246123 2307
rect 247064 2075 247249 2307
rect 247747 2075 247922 2307
rect 12943 1674 13184 1912
rect 248380 1343 248635 1577
rect 46480 677 46549 1236
rect 13322 -1699 46303 -1615
rect 46720 -1699 247871 -1615
rect 248379 -1715 248634 -1481
rect 248833 -1696 248940 -54
rect 12944 -2111 13185 -1873
rect 13323 -1976 46304 -1892
rect 46721 -1974 247872 -1890
rect -860 -5294 -704 -3774
rect 46474 -4774 46562 -4207
rect 12944 -5107 13185 -4869
rect 12944 -5504 13070 -5316
rect 23221 -5504 23406 -5316
rect 69528 -5504 69713 -5316
rect 122021 -5504 122206 -5316
rect 174621 -5504 174806 -5316
rect 230729 -5504 230914 -5316
rect 247793 -5504 247910 -5316
rect 13541 -5760 13741 -5572
rect 24116 -5760 24443 -5572
rect 70423 -5760 70750 -5572
rect 122916 -5760 123243 -5572
rect 175516 -5760 175843 -5572
rect 231624 -5760 231951 -5572
rect 247405 -5760 247587 -5572
<< metal3 >>
rect 13467 2614 13696 2928
rect 13467 2382 13479 2614
rect 13685 2382 13696 2614
rect 13467 2369 13696 2382
rect 13803 2307 14032 2928
rect 46289 2614 46871 2622
rect 46289 2382 46295 2614
rect 46381 2382 46777 2614
rect 46863 2382 46871 2614
rect 46289 2377 46871 2382
rect 13803 2075 13815 2307
rect 14021 2075 14032 2307
rect 13803 2059 14032 2075
rect 46288 2307 46872 2315
rect 46288 2075 46297 2307
rect 46383 2075 46777 2307
rect 46863 2075 46872 2307
rect 46288 2065 46872 2075
rect 53669 2307 53890 3112
rect 54547 2614 54910 3112
rect 54547 2382 54573 2614
rect 54892 2382 54910 2614
rect 54547 2361 54910 2382
rect 53669 2075 53688 2307
rect 53871 2075 53890 2307
rect 53669 2037 53890 2075
rect 164047 2307 164268 3112
rect 164942 2614 165304 3112
rect 164942 2382 164959 2614
rect 165286 2382 165304 2614
rect 164942 2361 165304 2382
rect 164047 2075 164064 2307
rect 164249 2075 164268 2307
rect 164047 2037 164268 2075
rect 231215 2307 231436 3113
rect 232110 2614 232472 3112
rect 232110 2382 232127 2614
rect 232454 2382 232472 2614
rect 232110 2361 232472 2382
rect 231215 2075 231232 2307
rect 231417 2075 231436 2307
rect 231215 2037 231436 2075
rect 236475 2307 236696 3112
rect 237370 2614 237728 3112
rect 237370 2382 237387 2614
rect 237714 2382 237728 2614
rect 237370 2361 237728 2382
rect 236475 2075 236492 2307
rect 236677 2075 236696 2307
rect 236475 2037 236696 2075
rect 239645 2307 239866 3112
rect 240540 2614 240898 3112
rect 240540 2382 240557 2614
rect 240884 2382 240898 2614
rect 240540 2361 240898 2382
rect 239645 2075 239662 2307
rect 239847 2075 239866 2307
rect 239645 2037 239866 2075
rect 241737 2307 241958 3112
rect 242632 2614 242990 3112
rect 242632 2382 242649 2614
rect 242976 2382 242990 2614
rect 242632 2361 242990 2382
rect 241737 2075 241754 2307
rect 241939 2075 241958 2307
rect 241737 2037 241958 2075
rect 243829 2307 244050 3112
rect 244724 2614 245082 3112
rect 244724 2382 244741 2614
rect 245068 2382 245082 2614
rect 244724 2361 245082 2382
rect 243829 2075 243846 2307
rect 244031 2075 244050 2307
rect 243829 2037 244050 2075
rect 245921 2307 246142 3112
rect 246276 2614 246634 3112
rect 246276 2382 246293 2614
rect 246620 2382 246634 2614
rect 246276 2361 246634 2382
rect 246705 2614 246944 3112
rect 246705 2382 246722 2614
rect 246894 2382 246944 2614
rect 246705 2361 246944 2382
rect 245921 2075 245938 2307
rect 246123 2075 246142 2307
rect 245921 2037 246142 2075
rect 247047 2307 247268 3112
rect 247389 2614 247632 3113
rect 247389 2382 247403 2614
rect 247620 2382 247632 2614
rect 247389 2362 247632 2382
rect 247047 2075 247064 2307
rect 247249 2075 247268 2307
rect 247047 2037 247268 2075
rect 247736 2307 247935 3114
rect 247736 2075 247747 2307
rect 247922 2075 247935 2307
rect 247736 2055 247935 2075
rect 12933 1912 13195 1940
rect 12933 1674 12943 1912
rect 13184 1674 13195 1912
rect 12933 -1873 13195 1674
rect 248367 1577 248645 1614
rect 248367 1343 248380 1577
rect 248635 1343 248645 1577
rect 46468 1236 46567 1304
rect 46468 677 46480 1236
rect 46549 677 46567 1236
rect 13297 -1526 46376 -1481
rect 13297 -1699 13322 -1526
rect 46303 -1699 46376 -1526
rect 13297 -1715 46376 -1699
rect 12933 -2111 12944 -1873
rect 13185 -1892 46376 -1873
rect 13185 -2065 13279 -1892
rect 46304 -2065 46376 -1892
rect 13185 -2111 46376 -2065
rect -1127 -3774 -681 -3754
rect -1127 -5294 -860 -3774
rect -704 -5294 -681 -3774
rect 12933 -4869 13195 -2111
rect 46468 -4207 46567 677
rect 248367 -1481 248645 1343
rect 46655 -1526 248379 -1481
rect 46655 -1700 46720 -1526
rect 247872 -1700 248379 -1526
rect 46655 -1715 248379 -1700
rect 248634 -1715 248645 -1481
rect 248804 -54 248973 -32
rect 248804 -1696 248833 -54
rect 248940 -1696 248973 -54
rect 248804 -1715 248973 -1696
rect 46655 -1889 248264 -1873
rect 46655 -2063 46720 -1889
rect 247872 -2063 248264 -1889
rect 46655 -2111 248264 -2063
rect 46468 -4774 46474 -4207
rect 46562 -4774 46567 -4207
rect 46468 -4780 46567 -4774
rect 12933 -5107 12944 -4869
rect 13185 -5107 13195 -4869
rect 248367 -5099 248645 -1715
rect 12933 -5141 13195 -5107
rect -1127 -5313 -681 -5294
rect 12937 -5316 13077 -5308
rect 12937 -5504 12944 -5316
rect 13070 -5504 13077 -5316
rect 12937 -5776 13077 -5504
rect 23204 -5316 23425 -5278
rect 23204 -5504 23221 -5316
rect 23406 -5504 23425 -5316
rect 13534 -5572 13749 -5550
rect 13534 -5760 13541 -5572
rect 13741 -5760 13749 -5572
rect 13534 -5935 13749 -5760
rect 23204 -6353 23425 -5504
rect 69511 -5316 69732 -5278
rect 69511 -5504 69528 -5316
rect 69713 -5504 69732 -5316
rect 24099 -5572 24461 -5551
rect 24099 -5760 24116 -5572
rect 24443 -5760 24461 -5572
rect 24099 -6353 24461 -5760
rect 69511 -6353 69732 -5504
rect 122004 -5316 122225 -5277
rect 122004 -5504 122021 -5316
rect 122206 -5504 122225 -5316
rect 70406 -5572 70768 -5551
rect 70406 -5760 70423 -5572
rect 70750 -5760 70768 -5572
rect 70406 -6353 70768 -5760
rect 122004 -6352 122225 -5504
rect 174604 -5316 174825 -5277
rect 174604 -5504 174621 -5316
rect 174806 -5504 174825 -5316
rect 122899 -5572 123261 -5550
rect 122899 -5760 122916 -5572
rect 123243 -5760 123261 -5572
rect 122899 -6352 123261 -5760
rect 174604 -6352 174825 -5504
rect 230712 -5316 230933 -5277
rect 230712 -5504 230729 -5316
rect 230914 -5504 230933 -5316
rect 175499 -5572 175861 -5550
rect 175499 -5760 175516 -5572
rect 175843 -5760 175861 -5572
rect 175499 -6352 175861 -5760
rect 230712 -6352 230933 -5504
rect 247785 -5316 247919 -5300
rect 247785 -5504 247793 -5316
rect 247910 -5504 247919 -5316
rect 231607 -5572 231969 -5550
rect 231607 -5760 231624 -5572
rect 231951 -5760 231969 -5572
rect 231607 -6352 231969 -5760
rect 247395 -5572 247600 -5553
rect 247395 -5760 247405 -5572
rect 247587 -5760 247600 -5572
rect 247395 -6160 247600 -5760
rect 247785 -6158 247919 -5504
<< via3 >>
rect 13322 -1615 46303 -1526
rect 13322 -1699 46303 -1615
rect 13279 -1976 13323 -1892
rect 13323 -1976 46304 -1892
rect 13279 -2065 46304 -1976
rect -860 -5294 -704 -3774
rect 46720 -1615 247872 -1526
rect 46720 -1699 247871 -1615
rect 247871 -1699 247872 -1615
rect 46720 -1700 247872 -1699
rect 248833 -1696 248940 -54
rect 46720 -1890 247872 -1889
rect 46720 -1974 46721 -1890
rect 46721 -1974 247872 -1890
rect 46720 -2063 247872 -1974
<< metal4 >>
rect -1132 -54 249191 -33
rect -1132 -1526 248833 -54
rect -1132 -1699 13322 -1526
rect 46303 -1699 46720 -1526
rect -1132 -1700 46720 -1699
rect 247872 -1696 248833 -1526
rect 248940 -1696 249191 -54
rect 247872 -1700 249191 -1696
rect -1132 -1718 249191 -1700
rect -1125 -1889 249191 -1869
rect -1125 -1892 46720 -1889
rect -1125 -2065 13279 -1892
rect 46304 -2063 46720 -1892
rect 247872 -2063 249191 -1889
rect 46304 -2065 249191 -2063
rect -1125 -3554 249191 -2065
rect -1127 -3774 -680 -3753
rect -1127 -5294 -860 -3774
rect -704 -5294 -680 -3774
rect -1127 -5313 -680 -5294
<< comment >>
rect 46354 -5615 46422 -5536
rect 46832 -5615 46900 -5536
rect 46354 -5773 46900 -5615
use bias_nstack  bias_nstack_0
array 0 439 -534 0 0 -3895
timestamp 1714090311
transform -1 0 17154 0 -1 -4733
box 3258 -2860 3926 1035
use bias_pstack  bias_pstack_0
array 0 439 534 0 0 -4355
timestamp 1714090311
transform 1 0 11201 0 -1 -1327
box 1986 -3967 2714 388
use sky130_fd_pr__res_high_po_0p35_P35QVK  XR2 paramcells
timestamp 1713888873
transform 1 0 6139 0 1 -1753
box -6758 -3582 6758 3582
<< labels >>
flabel metal3 164047 2871 164268 3112 0 FreeSans 1600 90 0 0 enb_10000_1
port 16 nsew
flabel metal3 164942 2871 165304 3112 0 FreeSans 1600 90 0 0 src_10000_1
port 15 nsew
flabel metal3 122004 -6352 122225 -6123 0 FreeSans 1600 90 0 0 ena_5000_1
port 33 nsew
flabel metal3 174604 -6352 174825 -6123 0 FreeSans 1600 90 0 0 ena_5000_2
port 35 nsew
flabel metal1 -902 1231 -702 1431 0 FreeSans 256 0 0 0 ref_in
port 1 nsew
flabel metal3 12937 -5776 13077 -5639 0 FreeSans 1600 90 0 0 ena_test0
port 39 nsew
flabel metal3 13534 -5935 13749 -5782 0 FreeSans 1600 90 0 0 snk_test0
port 40 nsew
flabel metal3 13467 2695 13696 2928 0 FreeSans 1600 90 0 0 src_test0
port 45 nsew
flabel metal3 13803 2695 14032 2928 0 FreeSans 1600 90 0 0 enb_test0
port 46 nsew
flabel metal3 122899 -6352 123261 -6123 0 FreeSans 1600 90 0 0 snk_5000_1
port 34 nsew
flabel metal3 175499 -6352 175861 -6123 0 FreeSans 1600 90 0 0 snk_5000_2
port 36 nsew
flabel metal3 23204 -6353 23425 -6124 0 FreeSans 1600 90 0 0 ena_2000
port 49 nsew
flabel metal3 24099 -6353 24461 -6124 0 FreeSans 1600 90 0 0 snk_2000
port 32 nsew
flabel metal2 35472 -5790 35672 -5590 0 FreeSans 256 0 0 0 ena
port 11 nsew
flabel metal2 46562 2684 46722 2884 0 FreeSans 256 0 0 0 enb
port 3 nsew
flabel comment 46623 -5695 46623 -5695 0 FreeSans 1600 0 0 0 mirror
flabel metal3 54548 2871 54910 3112 0 FreeSans 1600 90 0 0 src_10000_0
port 14 nsew
flabel metal3 53669 2897 53890 3112 0 FreeSans 1600 90 0 0 enb_10000_0
port 13 nsew
flabel metal3 69511 -6353 69732 -6124 0 FreeSans 1600 90 0 0 ena_5000_0
port 31 nsew
flabel metal3 70406 -6353 70768 -6124 0 FreeSans 1600 90 0 0 snk_5000_0
port 48 nsew
flabel metal3 231215 2872 231436 3113 0 FreeSans 1600 90 0 0 enb_600
port 17 nsew
flabel metal3 232110 2871 232472 3112 0 FreeSans 1600 90 0 0 src_600
port 18 nsew
flabel metal3 236475 2872 236696 3112 0 FreeSans 1600 90 0 0 enb_400
port 19 nsew
flabel metal3 237370 2872 237728 3112 0 FreeSans 1600 90 0 0 src_400
port 20 nsew
flabel metal3 239645 2872 239866 3112 0 FreeSans 1600 90 0 0 enb_200_0
port 21 nsew
flabel metal3 240540 2872 240898 3112 0 FreeSans 1600 90 0 0 src_200_0
port 22 nsew
flabel metal3 241737 2872 241958 3112 0 FreeSans 1600 90 0 0 enb_200_1
port 23 nsew
flabel metal3 242632 2872 242990 3112 0 FreeSans 1600 90 0 0 src_200_1
port 24 nsew
flabel metal3 243829 2872 244050 3112 0 FreeSans 1600 90 0 0 enb_200_2
port 25 nsew
flabel metal3 244724 2872 245082 3112 0 FreeSans 1600 90 0 0 src_200_2
port 26 nsew
flabel metal3 245921 2872 246142 3112 0 FreeSans 1600 90 0 0 enb_100
port 27 nsew
flabel metal3 246276 2872 246634 3112 0 FreeSans 1600 90 0 0 src_100
port 28 nsew
flabel metal3 246705 2872 246944 3112 0 FreeSans 1600 90 0 0 src_50
port 30 nsew
flabel metal3 247047 2872 247268 3112 0 FreeSans 1600 90 0 0 enb_50
port 29 nsew
flabel metal3 247736 2873 247935 3114 0 FreeSans 1600 90 0 0 enb_test1
port 44 nsew
flabel metal3 247389 2872 247632 3113 0 FreeSans 1600 90 0 0 src_test1
port 43 nsew
flabel metal3 247395 -6160 247600 -6018 0 FreeSans 1600 90 0 0 snk_test1
port 41 nsew
flabel metal3 247785 -6158 247919 -6016 0 FreeSans 1600 90 0 0 ena_test1
port 42 nsew
flabel metal3 230712 -6352 230933 -6164 0 FreeSans 1600 90 0 0 ena_3700
port 38 nsew
flabel metal3 231607 -6352 231969 -6164 0 FreeSans 1600 90 0 0 snk_3700
port 37 nsew
flabel metal4 -1132 -1718 -899 -33 0 FreeSans 1600 90 0 0 avdd
port 47 nsew
flabel metal4 -1125 -3554 -892 -1869 0 FreeSans 1600 90 0 0 avss
port 12 nsew
flabel metal4 -1127 -5313 -860 -3753 0 FreeSans 1600 90 0 0 vsub
port 50 nsew
<< end >>
