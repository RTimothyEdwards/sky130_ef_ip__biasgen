magic
tech sky130A
magscale 1 2
timestamp 1716925149
<< metal3 >>
rect -686 2492 686 2520
rect -686 1468 602 2492
rect 666 1468 686 2492
rect -686 1440 686 1468
rect -686 1172 686 1200
rect -686 148 602 1172
rect 666 148 686 1172
rect -686 120 686 148
rect -686 -148 686 -120
rect -686 -1172 602 -148
rect 666 -1172 686 -148
rect -686 -1200 686 -1172
rect -686 -1468 686 -1440
rect -686 -2492 602 -1468
rect 666 -2492 686 -1468
rect -686 -2520 686 -2492
<< via3 >>
rect 602 1468 666 2492
rect 602 148 666 1172
rect 602 -1172 666 -148
rect 602 -2492 666 -1468
<< mimcap >>
rect -646 2440 354 2480
rect -646 1520 -606 2440
rect 314 1520 354 2440
rect -646 1480 354 1520
rect -646 1120 354 1160
rect -646 200 -606 1120
rect 314 200 354 1120
rect -646 160 354 200
rect -646 -200 354 -160
rect -646 -1120 -606 -200
rect 314 -1120 354 -200
rect -646 -1160 354 -1120
rect -646 -1520 354 -1480
rect -646 -2440 -606 -1520
rect 314 -2440 354 -1520
rect -646 -2480 354 -2440
<< mimcapcontact >>
rect -606 1520 314 2440
rect -606 200 314 1120
rect -606 -1120 314 -200
rect -606 -2440 314 -1520
<< metal4 >>
rect -198 2441 -94 2640
rect 582 2492 686 2640
rect -607 2440 315 2441
rect -607 1520 -606 2440
rect 314 1520 315 2440
rect -607 1519 315 1520
rect -198 1121 -94 1519
rect 582 1468 602 2492
rect 666 1468 686 2492
rect 582 1172 686 1468
rect -607 1120 315 1121
rect -607 200 -606 1120
rect 314 200 315 1120
rect -607 199 315 200
rect -198 -199 -94 199
rect 582 148 602 1172
rect 666 148 686 1172
rect 582 -148 686 148
rect -607 -200 315 -199
rect -607 -1120 -606 -200
rect 314 -1120 315 -200
rect -607 -1121 315 -1120
rect -198 -1519 -94 -1121
rect 582 -1172 602 -148
rect 666 -1172 686 -148
rect 582 -1468 686 -1172
rect -607 -1520 315 -1519
rect -607 -2440 -606 -1520
rect 314 -2440 315 -1520
rect -607 -2441 315 -2440
rect -198 -2640 -94 -2441
rect 582 -2492 602 -1468
rect 666 -2492 686 -1468
rect 582 -2640 686 -2492
<< properties >>
string FIXED_BBOX -686 1440 394 2520
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 5.00 l 5.00 val 53.8 carea 2.00 cperi 0.19 nx 1 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
