magic
tech sky130A
magscale 1 2
timestamp 1719539418
<< error_s >>
rect 135078 -10275 135978 -9375
<< dnwell >>
rect 96152 17119 138230 24971
rect 89743 7919 138229 15771
rect 89743 -1281 138229 6571
rect 135078 -10481 138229 -2629
<< nwell >>
rect 96043 24765 138339 25080
rect 96043 17325 96358 24765
rect 138024 17325 138339 24765
rect 96043 17010 138339 17325
rect 89634 15565 138338 15880
rect 89634 8125 89949 15565
rect 138023 8125 138338 15565
rect 89634 7810 138338 8125
rect 89634 6365 138338 6680
rect 89634 -1075 89949 6365
rect 138023 -1075 138338 6365
rect 89634 -1390 138338 -1075
rect 135078 -2835 138338 -2520
rect 138023 -10275 138338 -2835
rect 135078 -10590 138338 -10275
<< pwell >>
rect 125398 17325 125486 17347
rect 108895 8125 108983 8147
rect 108895 -1075 108983 -1053
<< mvpsubdiff >>
rect 95923 25170 95983 25204
rect 137413 25170 137603 25204
rect 138399 25170 138459 25204
rect 95923 25144 95957 25170
rect 88137 24582 88197 24616
rect 95249 24582 95309 24616
rect 88137 24556 88171 24582
rect 88137 17652 88171 17678
rect 95275 24556 95309 24582
rect 95275 17652 95309 17678
rect 88137 17618 88197 17652
rect 95249 17618 95309 17652
rect 138425 25144 138459 25170
rect 95923 16898 95957 16924
rect 138425 16898 138459 16924
rect 95923 16864 95983 16898
rect 137413 16864 137603 16898
rect 138399 16864 138459 16898
rect 89514 15970 89574 16004
rect 90370 15970 90560 16004
rect 138398 15970 138458 16004
rect 89514 15944 89548 15970
rect 138424 15944 138458 15970
rect 89514 7698 89548 7724
rect 138424 7698 138458 7724
rect 89514 7664 89574 7698
rect 90370 7664 90560 7698
rect 138398 7664 138458 7698
rect 89514 6770 89574 6804
rect 90370 6770 90560 6804
rect 138398 6770 138458 6804
rect 89514 6744 89548 6770
rect 138424 6744 138458 6770
rect 89514 -1502 89548 -1476
rect 138424 -1502 138458 -1476
rect 89514 -1536 89574 -1502
rect 90370 -1536 90560 -1502
rect 138398 -1536 138458 -1502
rect 135144 -2430 135416 -2396
rect 138398 -2430 138458 -2396
rect 138424 -2456 138458 -2430
rect 138424 -10702 138458 -10676
rect 135144 -10736 135416 -10702
rect 138398 -10736 138458 -10702
<< mvnsubdiff >>
rect 96109 24994 138273 25014
rect 96109 24960 96189 24994
rect 137413 24960 137603 24994
rect 138193 24960 138273 24994
rect 96109 24940 138273 24960
rect 96109 24934 96183 24940
rect 96109 17156 96129 24934
rect 96163 17156 96183 24934
rect 96109 17150 96183 17156
rect 138199 24934 138273 24940
rect 138199 17156 138219 24934
rect 138253 17156 138273 24934
rect 138199 17150 138273 17156
rect 96109 17130 138273 17150
rect 96109 17096 96189 17130
rect 137413 17096 137603 17130
rect 138193 17096 138273 17130
rect 96109 17076 138273 17096
rect 89700 15794 138272 15814
rect 89700 15760 89780 15794
rect 90370 15760 90560 15794
rect 138192 15760 138272 15794
rect 89700 15740 138272 15760
rect 89700 15734 89774 15740
rect 89700 7956 89720 15734
rect 89754 7956 89774 15734
rect 89700 7950 89774 7956
rect 138198 15734 138272 15740
rect 138198 7956 138218 15734
rect 138252 7956 138272 15734
rect 138198 7950 138272 7956
rect 89700 7930 138272 7950
rect 89700 7896 89780 7930
rect 90370 7896 90560 7930
rect 138192 7896 138272 7930
rect 89700 7876 138272 7896
rect 89700 6594 138272 6614
rect 89700 6560 89780 6594
rect 90370 6560 90560 6594
rect 138192 6560 138272 6594
rect 89700 6540 138272 6560
rect 89700 6534 89774 6540
rect 89700 -1244 89720 6534
rect 89754 -1244 89774 6534
rect 89700 -1250 89774 -1244
rect 138198 6534 138272 6540
rect 138198 -1244 138218 6534
rect 138252 -1244 138272 6534
rect 138198 -1250 138272 -1244
rect 89700 -1270 138272 -1250
rect 89700 -1304 89780 -1270
rect 90370 -1304 90560 -1270
rect 138192 -1304 138272 -1270
rect 89700 -1324 138272 -1304
rect 135144 -2606 138272 -2586
rect 135144 -2640 135416 -2606
rect 138192 -2640 138272 -2606
rect 135144 -2660 138272 -2640
rect 138198 -2666 138272 -2660
rect 138198 -10444 138218 -2666
rect 138252 -10444 138272 -2666
rect 138198 -10450 138272 -10444
rect 135144 -10470 138272 -10450
rect 135144 -10504 135416 -10470
rect 138192 -10504 138272 -10470
rect 135144 -10524 138272 -10504
<< mvpsubdiffcont >>
rect 95983 25170 137413 25204
rect 137603 25170 138399 25204
rect 88197 24582 95249 24616
rect 88137 17678 88171 24556
rect 95275 17678 95309 24556
rect 88197 17618 95249 17652
rect 95923 16924 95957 25144
rect 138425 16924 138459 25144
rect 95983 16864 137413 16898
rect 137603 16864 138399 16898
rect 89574 15970 90370 16004
rect 90560 15970 138398 16004
rect 89514 7724 89548 15944
rect 138424 7724 138458 15944
rect 89574 7664 90370 7698
rect 90560 7664 138398 7698
rect 89574 6770 90370 6804
rect 90560 6770 138398 6804
rect 89514 -1476 89548 6744
rect 138424 -1476 138458 6744
rect 89574 -1536 90370 -1502
rect 90560 -1536 138398 -1502
rect 135416 -2430 138398 -2396
rect 138424 -10676 138458 -2456
rect 135416 -10736 138398 -10702
<< mvnsubdiffcont >>
rect 96189 24960 137413 24994
rect 137603 24960 138193 24994
rect 96129 17156 96163 24934
rect 138219 17156 138253 24934
rect 96189 17096 137413 17130
rect 137603 17096 138193 17130
rect 89780 15760 90370 15794
rect 90560 15760 138192 15794
rect 89720 7956 89754 15734
rect 138218 7956 138252 15734
rect 89780 7896 90370 7930
rect 90560 7896 138192 7930
rect 89780 6560 90370 6594
rect 90560 6560 138192 6594
rect 89720 -1244 89754 6534
rect 138218 -1244 138252 6534
rect 89780 -1304 90370 -1270
rect 90560 -1304 138192 -1270
rect 135416 -2640 138192 -2606
rect 138218 -10444 138252 -2666
rect 135416 -10504 138192 -10470
<< locali >>
rect 95923 25170 95983 25204
rect 137413 25170 137603 25204
rect 138399 25170 138459 25204
rect 95923 25155 138459 25170
rect 95923 25144 95969 25155
rect 88137 24582 88197 24616
rect 95249 24582 95923 24616
rect 88137 24556 95923 24582
rect 88171 24494 95275 24556
rect 88171 17740 88265 24494
rect 91871 23994 91918 24060
rect 94444 23994 94545 24059
rect 91871 23888 91879 23928
rect 90110 23166 90280 23182
rect 90110 23064 90131 23166
rect 90264 23064 90280 23166
rect 90110 23048 90280 23064
rect 92702 23166 92872 23182
rect 92702 23064 92723 23166
rect 92856 23064 92872 23166
rect 92702 23048 92872 23064
rect 91871 22366 91918 22432
rect 94453 22369 94554 22434
rect 91871 22257 91879 22297
rect 90110 21538 90280 21554
rect 90110 21436 90131 21538
rect 90264 21436 90280 21538
rect 90110 21420 90280 21436
rect 92702 21538 92872 21554
rect 92702 21436 92723 21538
rect 92856 21436 92872 21538
rect 92702 21420 92872 21436
rect 91871 20738 91918 20804
rect 94444 20737 94545 20802
rect 90110 19910 90280 19926
rect 90110 19808 90131 19910
rect 90264 19808 90280 19910
rect 90110 19792 90280 19808
rect 92702 19910 92872 19926
rect 92702 19808 92723 19910
rect 92856 19808 92872 19910
rect 92702 19792 92872 19808
rect 91871 19110 91918 19176
rect 94456 19109 94557 19174
rect 90110 18282 90280 18298
rect 90110 18180 90131 18282
rect 90264 18180 90280 18282
rect 90110 18164 90280 18180
rect 92702 18282 92872 18298
rect 92702 18180 92723 18282
rect 92856 18180 92872 18282
rect 92702 18164 92872 18180
rect 95192 17740 95275 24494
rect 88171 17678 95275 17740
rect 95309 24419 95923 24556
rect 95309 17678 95923 17814
rect 88137 17652 95923 17678
rect 88137 17618 88197 17652
rect 95249 17618 95923 17652
rect 95220 17617 95923 17618
rect 95957 16924 95969 25144
rect 95923 16914 95969 16924
rect 96021 25071 138361 25155
rect 96021 17010 96065 25071
rect 96129 24960 96189 24994
rect 137413 24960 137603 24994
rect 138193 24960 138253 24994
rect 96129 24934 138253 24960
rect 96163 24929 138219 24934
rect 96163 17156 96194 24929
rect 96129 17152 96194 17156
rect 96253 24892 138129 24929
rect 96253 24826 96850 24892
rect 97000 24826 138129 24892
rect 96253 24775 138129 24826
rect 96253 17309 96300 24775
rect 138082 17309 138129 24775
rect 96253 17152 138129 17309
rect 138188 17156 138219 24929
rect 138188 17152 138253 17156
rect 96129 17130 138253 17152
rect 96129 17096 96189 17130
rect 137413 17096 137603 17130
rect 138193 17096 138253 17130
rect 138317 17010 138361 25071
rect 96021 16923 138361 17010
rect 96021 16914 96074 16923
rect 95923 16898 96074 16914
rect 95923 16864 95983 16898
rect 137413 16864 137603 16923
rect 138308 16914 138361 16923
rect 138413 25144 138459 25155
rect 138413 16924 138425 25144
rect 138459 24419 138541 24616
rect 138459 17617 138541 17814
rect 138413 16914 138459 16924
rect 138308 16898 138459 16914
rect 138399 16864 138459 16898
rect 89514 15970 89574 16004
rect 90370 15970 90560 16004
rect 138398 15970 138458 16004
rect 89514 15955 138458 15970
rect 89514 15944 89560 15955
rect 89432 15219 89514 15416
rect 89432 8417 89514 8614
rect 89548 7724 89560 15944
rect 89514 7714 89560 7724
rect 89612 15871 138360 15955
rect 89612 7810 89656 15871
rect 89720 15760 89780 15794
rect 90370 15760 90560 15794
rect 138192 15760 138252 15794
rect 89720 15734 138252 15760
rect 89754 15729 138218 15734
rect 89754 7956 89785 15729
rect 89720 7952 89785 7956
rect 89844 15692 138128 15729
rect 89844 15626 137381 15692
rect 137531 15626 138128 15692
rect 89844 15575 138128 15626
rect 89844 8109 89891 15575
rect 138081 8109 138128 15575
rect 89844 7952 138128 8109
rect 138187 7956 138218 15729
rect 138187 7952 138252 7956
rect 89720 7930 138252 7952
rect 89720 7896 89780 7930
rect 90370 7896 90560 7930
rect 138192 7896 138252 7930
rect 138316 7810 138360 15871
rect 89612 7723 138360 7810
rect 89612 7714 89665 7723
rect 89514 7698 89665 7714
rect 89514 7664 89574 7698
rect 90370 7664 90560 7723
rect 138307 7714 138360 7723
rect 138412 15944 138458 15955
rect 138412 7724 138424 15944
rect 138458 15219 138540 15416
rect 138458 8417 138540 8614
rect 138412 7714 138458 7724
rect 138307 7698 138458 7714
rect 138398 7664 138458 7698
rect 89514 6770 89574 6804
rect 90370 6770 90560 6804
rect 138398 6770 138458 6804
rect 89514 6755 138458 6770
rect 89514 6744 89560 6755
rect 89432 6019 89514 6216
rect 89432 -783 89514 -586
rect 89548 -1476 89560 6744
rect 89514 -1486 89560 -1476
rect 89612 6671 138360 6755
rect 89612 -1390 89656 6671
rect 89720 6560 89780 6594
rect 90370 6560 90560 6594
rect 138192 6560 138252 6594
rect 89720 6534 138252 6560
rect 89754 6529 138218 6534
rect 89754 -1244 89785 6529
rect 89720 -1248 89785 -1244
rect 89844 6492 138128 6529
rect 89844 6426 137381 6492
rect 137531 6426 138128 6492
rect 89844 6375 138128 6426
rect 89844 -1091 89891 6375
rect 138081 -1091 138128 6375
rect 89844 -1248 138128 -1091
rect 138187 -1244 138218 6529
rect 138187 -1248 138252 -1244
rect 89720 -1270 138252 -1248
rect 89720 -1304 89780 -1270
rect 90370 -1304 90560 -1270
rect 138192 -1304 138252 -1270
rect 138316 -1390 138360 6671
rect 89612 -1477 138360 -1390
rect 89612 -1486 89665 -1477
rect 89514 -1502 89665 -1486
rect 89514 -1536 89574 -1502
rect 90370 -1536 90560 -1477
rect 138307 -1486 138360 -1477
rect 138412 6744 138458 6755
rect 138412 -1476 138424 6744
rect 138458 6019 138540 6216
rect 138458 -783 138540 -586
rect 138412 -1486 138458 -1476
rect 138307 -1502 138458 -1486
rect 138398 -1536 138458 -1502
rect 135144 -2430 135416 -2396
rect 138398 -2430 138458 -2396
rect 135144 -2445 138458 -2430
rect 135144 -2529 138360 -2445
rect 135152 -2640 135416 -2606
rect 138192 -2640 138252 -2606
rect 135152 -2666 138252 -2640
rect 135152 -2671 138218 -2666
rect 135152 -2825 138128 -2671
rect 138081 -10291 138128 -2825
rect 135144 -10448 138128 -10291
rect 138187 -10444 138218 -2671
rect 138187 -10448 138252 -10444
rect 135144 -10470 138252 -10448
rect 135144 -10504 135416 -10470
rect 138192 -10504 138252 -10470
rect 138316 -10590 138360 -2529
rect 135144 -10677 138360 -10590
rect 135144 -10736 135416 -10677
rect 138307 -10686 138360 -10677
rect 138412 -2456 138458 -2445
rect 138412 -10676 138424 -2456
rect 138458 -3181 138540 -2984
rect 138458 -9983 138540 -9786
rect 138412 -10686 138458 -10676
rect 138307 -10702 138458 -10686
rect 138398 -10736 138458 -10702
<< viali >>
rect 92206 24024 92252 24203
rect 94798 24024 94844 24203
rect 91823 23716 91871 23947
rect 94415 23716 94463 23947
rect 90131 23064 90264 23166
rect 92723 23064 92856 23166
rect 92206 22396 92252 22575
rect 94798 22396 94844 22575
rect 91823 22088 91871 22319
rect 94415 22088 94463 22319
rect 90131 21436 90264 21538
rect 92723 21436 92856 21538
rect 92206 20768 92252 20947
rect 94798 20768 94844 20947
rect 91823 20460 91871 20691
rect 94415 20460 94463 20691
rect 90131 19808 90264 19910
rect 92723 19808 92856 19910
rect 92206 19140 92252 19319
rect 94798 19140 94844 19319
rect 91823 18832 91871 19063
rect 94415 18832 94463 19063
rect 90131 18180 90264 18282
rect 92723 18180 92856 18282
rect 95969 16914 96021 25155
rect 96194 17152 96253 24929
rect 96850 24826 97000 24892
rect 138129 17152 138188 24929
rect 96074 16898 137413 16923
rect 96074 16879 137413 16898
rect 137603 16898 138308 16923
rect 138361 16914 138413 25155
rect 137603 16879 138308 16898
rect 89560 7714 89612 15955
rect 89785 7952 89844 15729
rect 137381 15626 137531 15692
rect 138128 7952 138187 15729
rect 89665 7698 90370 7723
rect 89665 7679 90370 7698
rect 90560 7698 138307 7723
rect 138360 7714 138412 15955
rect 90560 7679 138307 7698
rect 89560 -1486 89612 6755
rect 89785 -1248 89844 6529
rect 137381 6426 137531 6492
rect 138128 -1248 138187 6529
rect 89665 -1502 90370 -1477
rect 89665 -1521 90370 -1502
rect 90560 -1502 138307 -1477
rect 138360 -1486 138412 6755
rect 90560 -1521 138307 -1502
rect 138128 -10448 138187 -2671
rect 135416 -10702 138307 -10677
rect 138360 -10686 138412 -2445
rect 135416 -10721 138307 -10702
<< metal1 >>
rect 95933 25155 96049 25197
rect 88353 24431 95047 24445
rect 88353 24272 93083 24431
rect 94358 24272 95047 24431
rect 92201 24215 92265 24216
rect 92200 24214 92265 24215
rect 92200 24203 92207 24214
rect 92200 24024 92206 24203
rect 92200 24014 92207 24024
rect 92259 24014 92265 24214
rect 94789 24214 94853 24216
rect 93698 24065 94684 24116
rect 92200 24012 92259 24014
rect 91822 23953 91862 23960
rect 91807 23947 91883 23953
rect 91807 23716 91823 23947
rect 91871 23928 91883 23947
rect 92201 23929 92241 24012
rect 91871 23782 91947 23928
rect 93698 23782 93749 24065
rect 94414 23953 94454 23960
rect 94633 23957 94684 24065
rect 94789 24014 94795 24214
rect 94847 24014 94853 24214
rect 95287 24080 95299 24120
rect 94789 23993 94853 24014
rect 95293 23957 95299 24080
rect 91871 23731 93749 23782
rect 94399 23947 94475 23953
rect 91871 23728 91947 23731
rect 91871 23716 91883 23728
rect 91807 23710 91883 23716
rect 94399 23716 94415 23947
rect 94463 23824 94475 23947
rect 94633 23920 95299 23957
rect 95351 23920 95357 24120
rect 94633 23906 95310 23920
rect 94463 23784 95669 23824
rect 94463 23716 94475 23784
rect 94399 23710 94475 23716
rect 88364 23466 90501 23639
rect 91780 23466 95047 23639
rect 95663 23624 95669 23784
rect 95721 23624 95727 23824
rect 88811 23346 88829 23403
rect 89205 23346 95047 23403
rect 90110 23166 90280 23182
rect 90110 23064 90131 23166
rect 90264 23064 90280 23166
rect 90110 23048 90280 23064
rect 92702 23166 92872 23182
rect 92702 23064 92723 23166
rect 92856 23064 92872 23166
rect 92702 23048 92872 23064
rect 88364 22649 93085 22822
rect 94355 22649 95047 22822
rect 92199 22586 92265 22588
rect 94792 22586 94851 22587
rect 92199 22575 92207 22586
rect 92199 22396 92206 22575
rect 92199 22386 92207 22396
rect 92259 22386 92265 22586
rect 92200 22384 92259 22386
rect 91822 22325 91862 22330
rect 91807 22319 91883 22325
rect 91807 22088 91823 22319
rect 91871 22297 91883 22319
rect 92201 22301 92241 22384
rect 94098 22382 94586 22433
rect 94789 22396 94795 22586
rect 94847 22396 94853 22586
rect 95171 22448 95183 22488
rect 91871 22151 91947 22297
rect 94098 22151 94149 22382
rect 94414 22325 94454 22330
rect 91871 22100 94149 22151
rect 94399 22319 94475 22325
rect 91871 22097 91947 22100
rect 91871 22088 91883 22097
rect 91807 22082 91883 22088
rect 94399 22088 94415 22319
rect 94463 22196 94475 22319
rect 94535 22323 94586 22382
rect 94782 22386 94795 22396
rect 94847 22386 94855 22396
rect 94782 22356 94855 22386
rect 95177 22323 95183 22448
rect 94535 22288 95183 22323
rect 95235 22288 95241 22488
rect 94535 22272 95214 22288
rect 94463 22156 95563 22196
rect 94463 22088 94475 22156
rect 94399 22082 94475 22088
rect 88347 21838 90505 22011
rect 91784 21838 95047 22011
rect 95557 21996 95563 22156
rect 95615 21996 95621 22196
rect 88811 21718 88825 21775
rect 89205 21718 95047 21775
rect 90110 21538 90280 21554
rect 90110 21436 90131 21538
rect 90264 21436 90280 21538
rect 90110 21420 90280 21436
rect 92702 21538 92872 21554
rect 92702 21436 92723 21538
rect 92856 21436 92872 21538
rect 92702 21420 92872 21436
rect 88375 21022 93087 21195
rect 94357 21022 95047 21195
rect 92201 20959 92265 20960
rect 92200 20958 92265 20959
rect 94792 20958 94851 20959
rect 92200 20947 92207 20958
rect 92200 20768 92206 20947
rect 92259 20928 92265 20958
rect 92200 20758 92207 20768
rect 92259 20758 92265 20888
rect 94047 20764 94635 20815
rect 94789 20768 94795 20958
rect 94847 20789 94853 20958
rect 95048 20811 95060 20851
rect 92200 20756 92259 20758
rect 91822 20697 91862 20701
rect 91807 20691 91883 20697
rect 91807 20460 91823 20691
rect 91871 20658 91883 20691
rect 91871 20512 91939 20658
rect 94047 20512 94098 20764
rect 94414 20697 94454 20701
rect 91871 20461 94098 20512
rect 94399 20691 94475 20697
rect 91871 20460 91939 20461
rect 91807 20458 91939 20460
rect 94399 20460 94415 20691
rect 94463 20568 94475 20691
rect 94584 20687 94635 20764
rect 94782 20758 94795 20768
rect 94847 20758 94852 20789
rect 94782 20728 94852 20758
rect 95054 20687 95060 20811
rect 94584 20636 95060 20687
rect 95112 20651 95118 20851
rect 94463 20528 95481 20568
rect 94463 20460 94475 20528
rect 91807 20454 91883 20458
rect 94399 20454 94475 20460
rect 88358 20222 90501 20395
rect 91780 20222 95047 20395
rect 95475 20368 95481 20528
rect 95533 20368 95539 20568
rect 88811 20090 88822 20147
rect 89205 20090 95047 20147
rect 90110 19910 90280 19926
rect 90110 19808 90131 19910
rect 90264 19808 90280 19910
rect 90110 19792 90280 19808
rect 92702 19910 92872 19926
rect 92702 19808 92723 19910
rect 92856 19808 92872 19910
rect 92702 19792 92872 19808
rect 88391 19400 93083 19573
rect 94353 19400 95047 19573
rect 92199 19330 92265 19332
rect 94792 19330 94851 19331
rect 92199 19319 92207 19330
rect 92199 19140 92206 19319
rect 92259 19300 92265 19330
rect 92199 19130 92207 19140
rect 92259 19130 92265 19260
rect 93801 19161 94616 19212
rect 92200 19128 92259 19130
rect 91826 19069 91866 19076
rect 91810 19063 91883 19069
rect 91810 18832 91823 19063
rect 91871 19046 91883 19063
rect 91871 18901 91941 19046
rect 93801 18901 93852 19161
rect 94418 19069 94458 19076
rect 94565 19074 94616 19161
rect 94789 19130 94795 19330
rect 94847 19158 94853 19330
rect 94928 19185 94940 19225
rect 94847 19130 94852 19158
rect 94789 19114 94852 19130
rect 94934 19074 94940 19185
rect 91871 18850 93852 18901
rect 94402 19063 94475 19069
rect 91871 18846 91941 18850
rect 91871 18832 91883 18846
rect 91810 18826 91883 18832
rect 94402 18832 94415 19063
rect 94463 18940 94475 19063
rect 94565 19025 94940 19074
rect 94992 19025 94998 19225
rect 94565 19023 94956 19025
rect 94463 18900 95391 18940
rect 94463 18832 94475 18900
rect 94402 18826 94475 18832
rect 91787 18793 91890 18797
rect 88347 18583 90501 18756
rect 91780 18583 95047 18756
rect 95385 18740 95391 18900
rect 95443 18740 95449 18940
rect 95933 18912 95969 25155
rect 95759 18881 95969 18912
rect 88811 18462 88822 18519
rect 89205 18462 95047 18519
rect 90110 18282 90280 18298
rect 90110 18180 90131 18282
rect 90264 18180 90280 18282
rect 90110 18164 90280 18180
rect 92702 18282 92872 18298
rect 92702 18180 92723 18282
rect 92856 18180 92872 18282
rect 92702 18164 92872 18180
rect 88425 17861 93088 17939
rect 94360 17861 95047 17939
rect 95759 17742 95788 18881
rect 95759 17710 95969 17742
rect 95933 16914 95969 17710
rect 96021 16942 96049 25155
rect 138333 25155 138449 25197
rect 96150 24929 96288 24980
rect 96150 22699 96194 24929
rect 96253 22699 96288 24929
rect 138094 24929 138232 24980
rect 96837 24892 97016 24904
rect 96837 24826 96850 24892
rect 97000 24881 97016 24892
rect 97000 24829 97151 24881
rect 97000 24826 97016 24829
rect 96837 24816 97016 24826
rect 96150 21057 96166 22699
rect 96273 21057 96288 22699
rect 96150 17152 96194 21057
rect 96253 17152 96288 21057
rect 138094 22699 138129 24929
rect 138188 22699 138232 24929
rect 138094 21057 138109 22699
rect 138216 21057 138232 22699
rect 96150 17105 96288 17152
rect 97096 16942 97150 17246
rect 138094 17152 138129 21057
rect 138188 17152 138232 21057
rect 138094 17105 138232 17152
rect 138333 16942 138361 25155
rect 138413 18912 138449 25155
rect 138413 18881 138541 18912
rect 96021 16923 138361 16942
rect 96021 16914 96074 16923
rect 95933 16879 96074 16914
rect 137413 16879 137603 16923
rect 138308 16914 138361 16923
rect 138413 17710 138541 17742
rect 138413 16914 138449 17710
rect 138308 16879 138449 16914
rect 95933 16864 138449 16879
rect 89524 15955 89640 15997
rect 89524 9712 89560 15955
rect 89432 9681 89560 9712
rect 89432 8510 89560 8542
rect 89524 7714 89560 8510
rect 89612 7742 89640 15955
rect 138332 15955 138448 15997
rect 89741 15729 89879 15780
rect 89741 13499 89785 15729
rect 89844 13499 89879 15729
rect 138093 15729 138231 15780
rect 137365 15692 137544 15704
rect 137365 15681 137381 15692
rect 137230 15629 137381 15681
rect 137365 15626 137381 15629
rect 137531 15626 137544 15692
rect 137365 15616 137544 15626
rect 89741 11857 89757 13499
rect 89864 11857 89879 13499
rect 89741 7952 89785 11857
rect 89844 7952 89879 11857
rect 138093 13499 138128 15729
rect 138187 13499 138231 15729
rect 138093 11857 138108 13499
rect 138215 11857 138231 13499
rect 89741 7905 89879 7952
rect 137231 7742 137285 8046
rect 138093 7952 138128 11857
rect 138187 7952 138231 11857
rect 138093 7905 138231 7952
rect 138332 7742 138360 15955
rect 138412 9712 138448 15955
rect 138412 9681 138540 9712
rect 89612 7723 138360 7742
rect 89612 7714 89665 7723
rect 89524 7679 89665 7714
rect 90370 7679 90560 7723
rect 138307 7714 138360 7723
rect 138412 8510 138540 8542
rect 138412 7714 138448 8510
rect 138307 7679 138448 7714
rect 89524 7664 138448 7679
rect 89524 6755 89640 6797
rect 89524 512 89560 6755
rect 89432 481 89560 512
rect 89432 -690 89560 -658
rect 89524 -1486 89560 -690
rect 89612 -1458 89640 6755
rect 138332 6755 138448 6797
rect 89741 6529 89879 6580
rect 89741 4299 89785 6529
rect 89844 4299 89879 6529
rect 138093 6529 138231 6580
rect 137365 6492 137544 6504
rect 137365 6481 137381 6492
rect 137230 6429 137381 6481
rect 137365 6426 137381 6429
rect 137531 6426 137544 6492
rect 137365 6416 137544 6426
rect 89741 2657 89757 4299
rect 89864 2657 89879 4299
rect 89741 -1248 89785 2657
rect 89844 -1248 89879 2657
rect 138093 4299 138128 6529
rect 138187 4299 138231 6529
rect 138093 2657 138108 4299
rect 138215 2657 138231 4299
rect 89741 -1295 89879 -1248
rect 137231 -1458 137285 -1154
rect 138093 -1248 138128 2657
rect 138187 -1248 138231 2657
rect 138093 -1295 138231 -1248
rect 138332 -1458 138360 6755
rect 138412 512 138448 6755
rect 138412 481 138540 512
rect 89612 -1477 138360 -1458
rect 89612 -1486 89665 -1477
rect 89524 -1521 89665 -1486
rect 90370 -1521 90560 -1477
rect 138307 -1486 138360 -1477
rect 138412 -690 138540 -658
rect 138412 -1486 138448 -690
rect 138307 -1521 138448 -1486
rect 89524 -1536 138448 -1521
rect 138332 -2445 138448 -2403
rect 138093 -2671 138231 -2620
rect 138093 -4901 138128 -2671
rect 138187 -4901 138231 -2671
rect 138093 -6543 138108 -4901
rect 138215 -6543 138231 -4901
rect 138093 -10448 138128 -6543
rect 138187 -10448 138231 -6543
rect 138093 -10495 138231 -10448
rect 138332 -10658 138360 -2445
rect 138412 -8688 138448 -2445
rect 138412 -8719 138540 -8688
rect 135144 -10677 138360 -10658
rect 135144 -10721 135416 -10677
rect 138307 -10686 138360 -10677
rect 138412 -9890 138540 -9858
rect 138412 -10686 138448 -9890
rect 138307 -10721 138448 -10686
rect 135144 -10736 138448 -10721
<< via1 >>
rect 93083 24268 94358 24431
rect 92207 24203 92259 24214
rect 92207 24024 92252 24203
rect 92252 24024 92259 24203
rect 92207 24014 92259 24024
rect 94795 24203 94847 24214
rect 94795 24024 94798 24203
rect 94798 24024 94844 24203
rect 94844 24024 94847 24203
rect 94795 24014 94847 24024
rect 95299 23920 95351 24120
rect 90501 23447 91780 23664
rect 95669 23624 95721 23824
rect 88829 23346 89205 23403
rect 90131 23064 90264 23166
rect 92723 23064 92856 23166
rect 93085 22629 94355 22844
rect 92207 22575 92259 22586
rect 92207 22396 92252 22575
rect 92252 22396 92259 22575
rect 92207 22386 92259 22396
rect 94795 22575 94847 22586
rect 94795 22396 94798 22575
rect 94798 22396 94844 22575
rect 94844 22396 94847 22575
rect 94795 22386 94847 22396
rect 95183 22288 95235 22488
rect 90505 21820 91784 22037
rect 95563 21996 95615 22196
rect 88825 21718 89205 21775
rect 90131 21436 90264 21538
rect 92723 21436 92856 21538
rect 93087 21009 94357 21224
rect 92207 20947 92259 20958
rect 92207 20768 92252 20947
rect 92252 20768 92259 20947
rect 92207 20758 92259 20768
rect 94795 20947 94847 20958
rect 94795 20768 94798 20947
rect 94798 20768 94844 20947
rect 94844 20768 94847 20947
rect 94795 20758 94847 20768
rect 95060 20651 95112 20851
rect 90501 20189 91780 20406
rect 95481 20368 95533 20568
rect 88822 20090 89205 20147
rect 90131 19808 90264 19910
rect 92723 19808 92856 19910
rect 93083 19376 94353 19591
rect 92207 19319 92259 19330
rect 92207 19140 92252 19319
rect 92252 19140 92259 19319
rect 92207 19130 92259 19140
rect 94795 19319 94847 19330
rect 94795 19140 94798 19319
rect 94798 19140 94844 19319
rect 94844 19140 94847 19319
rect 94795 19130 94847 19140
rect 94940 19025 94992 19225
rect 90501 18563 91780 18780
rect 95391 18740 95443 18940
rect 88822 18462 89205 18519
rect 90131 18180 90264 18282
rect 92723 18180 92856 18282
rect 93088 17848 94360 17963
rect 95788 17742 95969 18881
rect 95969 17742 96002 18881
rect 96166 21057 96194 22699
rect 96194 21057 96253 22699
rect 96253 21057 96273 22699
rect 138109 21057 138129 22699
rect 138129 21057 138188 22699
rect 138188 21057 138216 22699
rect 138380 17742 138413 18881
rect 138413 17742 138541 18881
rect 89432 8542 89560 9681
rect 89560 8542 89593 9681
rect 89757 11857 89785 13499
rect 89785 11857 89844 13499
rect 89844 11857 89864 13499
rect 138108 11857 138128 13499
rect 138128 11857 138187 13499
rect 138187 11857 138215 13499
rect 138379 8542 138412 9681
rect 138412 8542 138540 9681
rect 89432 -658 89560 481
rect 89560 -658 89593 481
rect 89757 2657 89785 4299
rect 89785 2657 89844 4299
rect 89844 2657 89864 4299
rect 138108 2657 138128 4299
rect 138128 2657 138187 4299
rect 138187 2657 138215 4299
rect 138379 -658 138412 481
rect 138412 -658 138540 481
rect 138108 -6543 138128 -4901
rect 138128 -6543 138187 -4901
rect 138187 -6543 138215 -4901
rect 138379 -9858 138412 -8719
rect 138412 -9858 138540 -8719
<< metal2 >>
rect 92213 26130 103505 26178
rect 88811 24251 89205 24494
rect 88811 23403 88842 24251
rect 89174 23403 89205 24251
rect 88811 23346 88829 23403
rect 88811 23113 88842 23346
rect 89174 23113 89205 23346
rect 90488 23664 91793 24501
rect 92213 24224 92253 26130
rect 92351 26034 103347 26082
rect 92207 24214 92259 24224
rect 92207 24006 92259 24014
rect 90488 23447 90501 23664
rect 91780 23447 91793 23664
rect 92351 23594 92391 26034
rect 90110 23166 90280 23182
rect 90110 23139 90131 23166
rect 88811 21775 89205 23113
rect 88811 21718 88825 21775
rect 88811 20147 89205 21718
rect 88811 20090 88822 20147
rect 88811 18519 89205 20090
rect 88811 18462 88822 18519
rect 88811 17701 89205 18462
rect 89750 23099 90131 23139
rect 89750 17078 89790 23099
rect 90110 23064 90131 23099
rect 90264 23064 90280 23166
rect 90110 23048 90280 23064
rect 90488 22680 91793 23447
rect 90488 22037 90532 22680
rect 91734 22037 91793 22680
rect 92213 23554 92391 23594
rect 92478 25938 101890 25986
rect 92213 22596 92253 23554
rect 92478 23428 92518 25938
rect 92343 23388 92518 23428
rect 92597 25842 101702 25890
rect 92207 22586 92259 22596
rect 92207 22378 92259 22386
rect 92343 22187 92383 23388
rect 92597 23275 92637 25842
rect 94481 25746 100302 25794
rect 90488 21820 90505 22037
rect 91784 21820 91793 22037
rect 90110 21538 90280 21554
rect 90110 21497 90131 21538
rect 89870 21457 90131 21497
rect 89870 17078 89910 21457
rect 90110 21436 90131 21457
rect 90264 21436 90280 21538
rect 90110 21420 90280 21436
rect 90488 21089 90532 21820
rect 91734 21089 91793 21820
rect 90488 20406 91793 21089
rect 92213 22147 92383 22187
rect 92453 23235 92637 23275
rect 93070 24431 94373 24486
rect 93070 24268 93083 24431
rect 94358 24268 94373 24431
rect 92213 20968 92253 22147
rect 92453 21841 92493 23235
rect 92702 23166 92872 23182
rect 92702 23139 92723 23166
rect 92324 21801 92493 21841
rect 92602 23099 92723 23139
rect 92207 20958 92259 20968
rect 92207 20750 92259 20758
rect 92324 20646 92364 21801
rect 92602 21614 92642 23099
rect 92702 23064 92723 23099
rect 92856 23064 92872 23166
rect 92702 23048 92872 23064
rect 90488 20189 90501 20406
rect 91780 20189 91793 20406
rect 90110 19910 90280 19926
rect 90110 19874 90131 19910
rect 89990 19834 90131 19874
rect 89990 17078 90030 19834
rect 90110 19808 90131 19834
rect 90264 19808 90280 19910
rect 90110 19792 90280 19808
rect 90488 18780 91793 20189
rect 92213 20606 92364 20646
rect 92482 21574 92642 21614
rect 93070 22844 94373 24268
rect 93070 22629 93085 22844
rect 94355 22629 94373 22844
rect 92213 19340 92253 20606
rect 92482 20166 92522 21574
rect 92702 21538 92872 21554
rect 92702 21497 92723 21538
rect 92342 20126 92522 20166
rect 92601 21457 92723 21497
rect 92207 19330 92259 19340
rect 92207 19122 92259 19130
rect 90488 18563 90501 18780
rect 91780 18563 91793 18780
rect 90110 18282 90280 18298
rect 90110 18180 90131 18282
rect 90264 18180 90280 18282
rect 90110 18164 90280 18180
rect 90110 17078 90150 18164
rect 90488 17790 91793 18563
rect 92342 17078 92382 20126
rect 92601 20045 92641 21457
rect 92702 21436 92723 21457
rect 92856 21436 92872 21538
rect 92702 21420 92872 21436
rect 92462 20005 92641 20045
rect 93070 21224 94373 22629
rect 93070 21009 93087 21224
rect 94357 21009 94373 21224
rect 92462 17078 92502 20005
rect 92702 19910 92872 19926
rect 92702 19874 92723 19910
rect 92578 19834 92723 19874
rect 92578 17496 92622 19834
rect 92702 19808 92723 19834
rect 92856 19808 92872 19910
rect 92702 19792 92872 19808
rect 93070 19591 94373 21009
rect 94481 20490 94521 25746
rect 94667 25650 100166 25698
rect 94667 22270 94707 25650
rect 94801 25554 98652 25602
rect 94801 24224 94841 25554
rect 94937 25458 98496 25506
rect 94795 24214 94847 24224
rect 94795 24006 94847 24014
rect 94937 23784 94977 25458
rect 97268 25135 97875 25367
rect 98178 25135 98400 25367
rect 97089 24828 97688 25060
rect 97832 25043 98400 25060
rect 98448 25043 98496 25458
rect 97832 24995 98496 25043
rect 98604 25060 98652 25554
rect 98813 25135 99452 25367
rect 99473 25134 100025 25367
rect 98604 25003 99348 25060
rect 97832 24828 98400 24995
rect 98663 24828 99348 25003
rect 99742 25044 99837 25060
rect 100118 25044 100166 25650
rect 99742 24996 100166 25044
rect 100254 25060 100302 25746
rect 100455 25135 101556 25367
rect 99742 24989 99837 24996
rect 99741 24828 99837 24989
rect 100254 24828 100920 25060
rect 101347 25049 101556 25060
rect 101654 25049 101702 25842
rect 101347 25001 101702 25049
rect 101842 25060 101890 25938
rect 102053 25135 103234 25367
rect 101347 24828 101556 25001
rect 101842 24984 102516 25060
rect 101882 24828 102516 24984
rect 102961 25040 103139 25060
rect 103299 25040 103347 26034
rect 102961 24992 103347 25040
rect 103457 25060 103505 26130
rect 103660 25135 130926 25367
rect 131253 25135 137417 25367
rect 102961 24828 103139 24992
rect 103457 24981 137257 25060
rect 103481 24828 137257 24981
rect 97847 24827 97887 24828
rect 100254 24827 100302 24828
rect 96765 24427 137661 24665
rect 95299 24120 95351 24128
rect 96442 24096 96471 24330
rect 96726 24096 96773 24330
rect 137539 24096 137661 24330
rect 137911 24096 137940 24330
rect 95299 23914 95351 23920
rect 95300 23907 95345 23914
rect 94937 23744 94979 23784
rect 94937 23578 94977 23744
rect 94801 23538 94977 23578
rect 94801 22596 94841 23538
rect 94795 22586 94847 22596
rect 94795 22378 94847 22386
rect 95183 22488 95235 22496
rect 95183 22282 95235 22288
rect 95184 22275 95229 22282
rect 94667 22230 94841 22270
rect 94801 20968 94841 22230
rect 94795 20958 94847 20968
rect 94795 20750 94847 20758
rect 95060 20851 95112 20859
rect 95058 20651 95060 20688
rect 95058 20645 95112 20651
rect 95058 20638 95106 20645
rect 94481 20450 94841 20490
rect 93070 19376 93083 19591
rect 94353 19376 94373 19591
rect 93070 18885 94373 19376
rect 94801 19340 94841 20450
rect 94795 19330 94847 19340
rect 94795 19122 94847 19130
rect 94940 19225 94992 19233
rect 94940 19019 94992 19025
rect 92702 18282 92872 18298
rect 92702 18180 92723 18282
rect 92856 18180 92872 18282
rect 92702 18164 92872 18180
rect 92578 17078 92618 17496
rect 92702 17078 92742 18164
rect 93070 17963 93104 18885
rect 94346 17963 94373 18885
rect 93070 17848 93088 17963
rect 94360 17848 94373 17963
rect 93070 17740 93104 17848
rect 94346 17740 94373 17848
rect 93070 17700 94373 17740
rect 94943 19012 94986 19019
rect 94943 16305 94982 19012
rect 95058 16400 95097 20638
rect 95184 16496 95223 22275
rect 95300 16592 95339 23907
rect 95669 23824 95721 23832
rect 95669 23618 95721 23624
rect 95563 22196 95615 22204
rect 95563 21990 95615 21996
rect 95481 20568 95533 20576
rect 95481 20362 95533 20368
rect 95391 18940 95443 18948
rect 95391 18734 95443 18740
rect 95397 16690 95437 18734
rect 95487 16780 95527 20362
rect 95569 16862 95609 21990
rect 95675 16948 95715 23618
rect 96765 23096 137661 23330
rect 137541 23095 137661 23096
rect 96111 22699 96302 22722
rect 96111 21057 96166 22699
rect 96273 21057 96302 22699
rect 138080 22699 138271 22722
rect 96765 22092 137617 22326
rect 96111 21038 96302 21057
rect 96443 21038 96472 21272
rect 96727 21038 96773 21272
rect 137545 21138 137655 21272
rect 137413 21054 137655 21138
rect 137545 21038 137655 21054
rect 137910 21038 137939 21272
rect 138080 21057 138109 22699
rect 138216 21057 138271 22699
rect 138080 21038 138271 21057
rect 126302 20863 137661 20880
rect 137413 20779 137661 20863
rect 137335 20777 137661 20779
rect 126302 20642 137661 20777
rect 96784 19618 137605 19856
rect 95759 18881 96023 18912
rect 95759 17742 95788 18881
rect 96002 17742 96023 18881
rect 138359 18881 138541 18912
rect 95759 17710 96023 17742
rect 96784 17646 137661 17884
rect 138359 17742 138380 18881
rect 138359 17710 138541 17742
rect 97081 17249 97691 17437
rect 98171 17379 98770 17437
rect 98152 17249 98770 17379
rect 99209 17317 99839 17437
rect 99201 17249 99839 17317
rect 100278 17249 100909 17437
rect 101348 17318 137222 17437
rect 101334 17249 137222 17318
rect 97246 16993 97856 17181
rect 98152 16948 98192 17249
rect 98300 16993 98935 17181
rect 95675 16908 98192 16948
rect 99201 16862 99241 17249
rect 99374 16993 99996 17181
rect 95569 16822 99241 16862
rect 100279 16780 100319 17249
rect 100435 16993 101072 17181
rect 95487 16740 100319 16780
rect 101334 16690 101374 17249
rect 132640 17181 132967 17187
rect 101511 16993 137385 17181
rect 95397 16650 101374 16690
rect 95300 16553 96005 16592
rect 95184 16457 96005 16496
rect 95058 16361 96005 16400
rect 94943 16266 96005 16305
rect 90556 15936 136203 16167
rect 90556 15935 103128 15936
rect 103455 15935 136203 15936
rect 136506 15935 137113 16167
rect 134356 15934 134908 15935
rect 90716 15628 136549 15860
rect 136693 15628 137292 15860
rect 136494 15627 136534 15628
rect 90312 15227 137616 15465
rect 90033 14896 90062 15130
rect 90317 14896 90434 15130
rect 137608 14896 137655 15130
rect 137910 14896 137939 15130
rect 90312 13896 137616 14130
rect 90312 13895 90432 13896
rect 89702 13499 89893 13522
rect 89702 11857 89757 13499
rect 89864 11857 89893 13499
rect 138079 13499 138270 13522
rect 90356 12892 137616 13126
rect 89702 11838 89893 11857
rect 90034 11838 90063 12072
rect 90318 11938 90364 12072
rect 90318 11854 90560 11938
rect 90318 11838 90364 11854
rect 137608 11838 137654 12072
rect 137909 11838 137938 12072
rect 138079 11857 138108 13499
rect 138215 11857 138270 13499
rect 138079 11838 138270 11857
rect 90312 11663 108079 11680
rect 90312 11579 90560 11663
rect 90312 11577 90638 11579
rect 90312 11442 108079 11577
rect 90368 10418 137597 10656
rect 89432 9681 89614 9712
rect 89593 8542 89614 9681
rect 138358 9681 138540 9712
rect 89432 8510 89614 8542
rect 90312 8446 137597 8684
rect 138358 8542 138379 9681
rect 138358 8510 138540 8542
rect 90751 8049 136222 8237
rect 136690 8049 137300 8237
rect 101414 7981 101741 7987
rect 90588 7793 136081 7981
rect 136525 7793 137135 7981
rect 90556 6735 137113 6967
rect 134356 6734 134908 6735
rect 90716 6428 137292 6660
rect 136494 6427 136534 6428
rect 90312 6027 137616 6265
rect 90033 5696 90062 5930
rect 90317 5696 90434 5930
rect 137608 5696 137655 5930
rect 137910 5696 137939 5930
rect 90312 4696 137616 4930
rect 90312 4695 90432 4696
rect 89702 4299 89893 4322
rect 89702 2657 89757 4299
rect 89864 2657 89893 4299
rect 138079 4299 138270 4322
rect 90356 3692 137616 3926
rect 89702 2638 89893 2657
rect 90034 2638 90063 2872
rect 90318 2738 90364 2872
rect 90318 2654 90560 2738
rect 90318 2638 90364 2654
rect 137608 2638 137654 2872
rect 137909 2638 137938 2872
rect 138079 2657 138108 4299
rect 138215 2657 138270 4299
rect 138079 2638 138270 2657
rect 90312 2463 108079 2480
rect 90312 2379 90560 2463
rect 90312 2377 90638 2379
rect 90312 2242 108079 2377
rect 90368 1218 137597 1456
rect 89432 481 89614 512
rect 89593 -658 89614 481
rect 138358 481 138540 512
rect 89432 -690 89614 -658
rect 90312 -754 137597 -516
rect 138358 -658 138379 481
rect 138358 -690 138540 -658
rect 90751 -1151 136216 -963
rect 136690 -1151 137300 -963
rect 101414 -1219 101741 -1213
rect 90588 -1407 136081 -1219
rect 136525 -1407 137135 -1219
rect 135412 -2465 137704 -2233
rect 135572 -2772 137704 -2540
rect 135168 -3173 137704 -2935
rect 135168 -3504 135290 -3270
rect 137608 -3504 137655 -3270
rect 137910 -3504 137939 -3270
rect 135168 -4504 137704 -4270
rect 135168 -4505 135288 -4504
rect 138079 -4901 138270 -4878
rect 135224 -5508 137704 -5274
rect 137608 -6462 137654 -6328
rect 135215 -6546 135416 -6462
rect 137608 -6562 137654 -6546
rect 137909 -6562 137938 -6328
rect 138079 -6543 138108 -4901
rect 138215 -6543 138270 -4901
rect 138079 -6562 138270 -6543
rect 135168 -6737 137704 -6720
rect 135168 -6821 135416 -6737
rect 135168 -6823 135494 -6821
rect 135168 -6958 137704 -6823
rect 135224 -7982 137704 -7744
rect 138358 -8719 138540 -8688
rect 135168 -9954 137704 -9716
rect 138358 -9858 138379 -8719
rect 138358 -9890 138540 -9858
rect 135607 -10351 137704 -10163
rect 135444 -10607 137704 -10419
<< via2 >>
rect 88842 23403 89174 24251
rect 88842 23346 89174 23403
rect 88842 23113 89174 23346
rect 90532 22037 91734 22680
rect 90532 21820 91734 22037
rect 90532 21089 91734 21820
rect 130926 25135 131253 25367
rect 96471 24096 96726 24330
rect 137661 24096 137911 24330
rect 93104 17963 94346 18885
rect 93104 17848 94346 17963
rect 93104 17740 94346 17848
rect 96166 21057 96273 22699
rect 96472 21038 96727 21272
rect 97235 21054 137413 21138
rect 137655 21038 137910 21272
rect 138109 21057 138216 22699
rect 97234 20779 137413 20863
rect 125319 20777 137335 20779
rect 95788 17742 96002 18881
rect 138380 17742 138541 18881
rect 90062 14896 90317 15130
rect 137655 14896 137910 15130
rect 89757 11857 89864 13499
rect 90063 11838 90318 12072
rect 90560 11854 137146 11938
rect 137654 11838 137909 12072
rect 138108 11857 138215 13499
rect 90560 11579 137147 11663
rect 90638 11577 109062 11579
rect 89432 8542 89593 9681
rect 138379 8542 138540 9681
rect 90062 5696 90317 5930
rect 137655 5696 137910 5930
rect 89757 2657 89864 4299
rect 90063 2638 90318 2872
rect 90560 2654 137146 2738
rect 137654 2638 137909 2872
rect 138108 2657 138215 4299
rect 90560 2379 137147 2463
rect 90638 2377 109062 2379
rect 89432 -658 89593 481
rect 138379 -658 138540 481
rect 137655 -3504 137910 -3270
rect 137654 -6462 137909 -6328
rect 135416 -6546 137909 -6462
rect 137654 -6562 137909 -6546
rect 138108 -6543 138215 -4901
rect 135416 -6821 137704 -6737
rect 135494 -6823 137704 -6821
rect 138379 -9858 138540 -8719
<< metal3 >>
rect 130911 25500 131271 25752
rect 130912 25367 131270 25500
rect 130912 25135 130926 25367
rect 131253 25135 131270 25367
rect 130912 25114 131270 25135
rect 96461 24330 96739 24367
rect 88812 24251 89205 24286
rect 88812 23113 88842 24251
rect 89174 23113 89205 24251
rect 88812 23084 89205 23113
rect 96461 24096 96471 24330
rect 96726 24096 96739 24330
rect 90487 22680 91793 22723
rect 90487 21089 90532 22680
rect 91734 21089 91793 22680
rect 90487 21036 91793 21089
rect 96133 22699 96302 22721
rect 96133 21057 96166 22699
rect 96273 21057 96302 22699
rect 96133 21038 96302 21057
rect 96461 21272 96739 24096
rect 137643 24330 137921 24367
rect 137643 24096 137661 24330
rect 137911 24096 137921 24330
rect 137643 21272 137921 24096
rect 96461 21038 96472 21272
rect 96727 21227 137655 21272
rect 96727 21053 97234 21227
rect 137413 21053 137655 21227
rect 96727 21038 137655 21053
rect 137910 21038 137921 21272
rect 138080 22699 138249 22721
rect 138080 21057 138109 22699
rect 138216 21057 138249 22699
rect 138080 21038 138249 21057
rect 93072 18885 94372 18913
rect 93072 17740 93104 18885
rect 94346 17740 94372 18885
rect 93072 17713 94372 17740
rect 95759 18881 96023 18912
rect 95759 17742 95788 18881
rect 96002 17742 96023 18881
rect 95759 17710 96023 17742
rect 96461 17654 96739 21038
rect 96842 20864 137538 20880
rect 96842 20690 97234 20864
rect 137413 20690 137538 20864
rect 96842 20688 125319 20690
rect 137335 20688 137538 20690
rect 96842 20642 137538 20688
rect 137643 17654 137921 21038
rect 138359 18881 138547 18912
rect 138359 17742 138380 18881
rect 138541 17742 138547 18881
rect 138359 17710 138547 17742
rect 90052 15130 90330 15167
rect 90052 14896 90062 15130
rect 90317 14896 90330 15130
rect 89724 13499 89893 13521
rect 89724 11857 89757 13499
rect 89864 11857 89893 13499
rect 89724 11838 89893 11857
rect 90052 12072 90330 14896
rect 137642 15130 137920 15167
rect 137642 14896 137655 15130
rect 137910 14896 137920 15130
rect 137642 12072 137920 14896
rect 90052 11838 90063 12072
rect 90318 12027 137654 12072
rect 90318 11853 90560 12027
rect 137147 11853 137654 12027
rect 90318 11838 137654 11853
rect 137909 11838 137920 12072
rect 138079 13499 138248 13521
rect 138079 11857 138108 13499
rect 138215 11857 138248 13499
rect 138079 11838 138248 11857
rect 89427 9681 89614 9712
rect 89427 8542 89432 9681
rect 89593 8542 89614 9681
rect 89427 8510 89614 8542
rect 90052 8454 90330 11838
rect 90406 11664 137539 11680
rect 90406 11490 90560 11664
rect 137147 11490 137539 11664
rect 90406 11488 90638 11490
rect 109062 11488 137539 11490
rect 90406 11442 137539 11488
rect 137642 8454 137920 11838
rect 138358 9681 138545 9712
rect 138358 8542 138379 9681
rect 138540 8542 138545 9681
rect 138358 8510 138545 8542
rect 90052 5930 90330 5967
rect 90052 5696 90062 5930
rect 90317 5696 90330 5930
rect 89724 4299 89893 4321
rect 89724 2657 89757 4299
rect 89864 2657 89893 4299
rect 89724 2638 89893 2657
rect 90052 2872 90330 5696
rect 137642 5930 137920 5967
rect 137642 5696 137655 5930
rect 137910 5696 137920 5930
rect 137642 2872 137920 5696
rect 90052 2638 90063 2872
rect 90318 2827 137654 2872
rect 90318 2653 90560 2827
rect 137147 2653 137654 2827
rect 90318 2638 137654 2653
rect 137909 2638 137920 2872
rect 138079 4299 138248 4321
rect 138079 2657 138108 4299
rect 138215 2657 138248 4299
rect 138079 2638 138248 2657
rect 89427 481 89614 512
rect 89427 -658 89432 481
rect 89593 -658 89614 481
rect 89427 -690 89614 -658
rect 90052 -746 90330 2638
rect 90417 2464 137539 2480
rect 90417 2290 90560 2464
rect 137147 2290 137539 2464
rect 90417 2288 90638 2290
rect 109062 2288 137539 2290
rect 90417 2242 137539 2288
rect 137642 -746 137920 2638
rect 138358 481 138545 512
rect 138358 -658 138379 481
rect 138540 -658 138545 481
rect 138358 -690 138545 -658
rect 137642 -3270 137920 -3233
rect 137642 -3504 137655 -3270
rect 137910 -3504 137920 -3270
rect 137642 -6328 137920 -3504
rect 135208 -6373 137654 -6328
rect 135208 -6547 135416 -6373
rect 135208 -6562 137654 -6547
rect 137909 -6562 137920 -6328
rect 138079 -4901 138248 -4879
rect 138079 -6543 138108 -4901
rect 138215 -6543 138248 -4901
rect 138079 -6562 138248 -6543
rect 137642 -6720 137920 -6562
rect 135219 -6736 137920 -6720
rect 135219 -6910 135416 -6736
rect 135219 -6912 135494 -6910
rect 137704 -6912 137920 -6736
rect 135219 -6958 137920 -6912
rect 137642 -9946 137920 -6958
rect 138358 -8719 138545 -8688
rect 138358 -9858 138379 -8719
rect 138540 -9858 138545 -8719
rect 138358 -9890 138545 -9858
<< via3 >>
rect 88842 23113 89174 24251
rect 90532 21089 91734 22680
rect 96166 21057 96273 22699
rect 97234 21138 137413 21227
rect 97234 21054 97235 21138
rect 97235 21054 137413 21138
rect 97234 21053 137413 21054
rect 138109 21057 138216 22699
rect 93104 17740 94346 18885
rect 95788 17742 96002 18881
rect 97234 20863 137413 20864
rect 97234 20779 137413 20863
rect 97234 20777 125319 20779
rect 125319 20777 137335 20779
rect 137335 20777 137413 20779
rect 97234 20690 137413 20777
rect 125319 20688 137335 20690
rect 138380 17742 138541 18881
rect 89757 11857 89864 13499
rect 90560 11938 137147 12027
rect 90560 11854 137146 11938
rect 137146 11854 137147 11938
rect 90560 11853 137147 11854
rect 138108 11857 138215 13499
rect 89432 8542 89593 9681
rect 90560 11663 137147 11664
rect 90560 11579 137147 11663
rect 90560 11577 90638 11579
rect 90638 11577 109062 11579
rect 109062 11577 137147 11579
rect 90560 11490 137147 11577
rect 90638 11488 109062 11490
rect 138379 8542 138540 9681
rect 89757 2657 89864 4299
rect 90560 2738 137147 2827
rect 90560 2654 137146 2738
rect 137146 2654 137147 2738
rect 90560 2653 137147 2654
rect 138108 2657 138215 4299
rect 89432 -658 89593 481
rect 90560 2463 137147 2464
rect 90560 2379 137147 2463
rect 90560 2377 90638 2379
rect 90638 2377 109062 2379
rect 109062 2377 137147 2379
rect 90560 2290 137147 2377
rect 90638 2288 109062 2290
rect 138379 -658 138540 481
rect 135416 -6462 137654 -6373
rect 137654 -6462 137704 -6373
rect 135416 -6546 137704 -6462
rect 135416 -6547 137654 -6546
rect 137654 -6547 137704 -6546
rect 138108 -6543 138215 -4901
rect 135416 -6737 137704 -6736
rect 135416 -6821 137704 -6737
rect 135416 -6823 135494 -6821
rect 135494 -6823 137704 -6821
rect 135416 -6910 137704 -6823
rect 135494 -6912 137704 -6910
rect 138379 -9858 138540 -8719
<< metal4 >>
rect 88136 24251 96025 24283
rect 88136 23113 88842 24251
rect 89174 23113 96025 24251
rect 88136 23083 96025 23113
rect 138357 23083 138541 24283
rect 88136 22699 138541 22720
rect 88136 22680 96166 22699
rect 88136 21089 90532 22680
rect 91734 21089 96166 22680
rect 88136 21057 96166 21089
rect 96273 21227 138109 22699
rect 96273 21057 97234 21227
rect 88136 21053 97234 21057
rect 137413 21057 138109 21227
rect 138216 21057 138541 22699
rect 137413 21053 138541 21057
rect 88136 21035 138541 21053
rect 88136 20864 138541 20884
rect 88136 20690 97234 20864
rect 137413 20690 138541 20864
rect 88136 20688 125319 20690
rect 137335 20688 138541 20690
rect 88136 19199 138541 20688
rect 88136 18885 96025 18911
rect 88136 17740 93104 18885
rect 94346 18881 96025 18885
rect 94346 17742 95788 18881
rect 96002 17742 96025 18881
rect 94346 17740 96025 17742
rect 88136 17711 96025 17740
rect 138357 18881 138545 18911
rect 138357 17742 138380 18881
rect 138541 17742 138545 18881
rect 138357 17711 138545 17742
rect 89432 13883 89616 15083
rect 138356 13883 138540 15083
rect 89432 13499 138540 13520
rect 89432 11857 89757 13499
rect 89864 12027 138108 13499
rect 89864 11857 90560 12027
rect 89432 11853 90560 11857
rect 137147 11857 138108 12027
rect 138215 11857 138540 13499
rect 137147 11853 138540 11857
rect 89432 11835 138540 11853
rect 89432 11664 138540 11684
rect 89432 11490 90560 11664
rect 137147 11490 138540 11664
rect 89432 11488 90638 11490
rect 109062 11488 138540 11490
rect 89432 9999 138540 11488
rect 89429 9681 89616 9711
rect 89429 8542 89432 9681
rect 89593 8542 89616 9681
rect 89429 8511 89616 8542
rect 138356 9681 138544 9711
rect 138356 8542 138379 9681
rect 138540 8542 138544 9681
rect 138356 8511 138544 8542
rect 89432 4683 89616 5883
rect 138356 4683 138540 5883
rect 89432 4299 138540 4320
rect 89432 2657 89757 4299
rect 89864 2827 138108 4299
rect 89864 2657 90560 2827
rect 89432 2653 90560 2657
rect 137147 2657 138108 2827
rect 138215 2657 138540 4299
rect 137147 2653 138540 2657
rect 89432 2635 138540 2653
rect 89432 2464 138540 2484
rect 89432 2290 90560 2464
rect 137147 2290 138540 2464
rect 89432 2288 90638 2290
rect 109062 2288 138540 2290
rect 89432 799 138540 2288
rect 89429 481 89616 511
rect 89429 -658 89432 481
rect 89593 -658 89616 481
rect 89429 -689 89616 -658
rect 138356 481 138543 511
rect 138356 -658 138379 481
rect 138540 -658 138543 481
rect 138356 -689 138543 -658
rect 138356 -4517 138540 -3317
rect 135167 -4901 138540 -4880
rect 135167 -6373 138108 -4901
rect 135167 -6547 135416 -6373
rect 137704 -6543 138108 -6373
rect 138215 -6543 138540 -4901
rect 137704 -6547 138540 -6543
rect 135167 -6565 138540 -6547
rect 135168 -6736 138540 -6716
rect 135168 -6910 135416 -6736
rect 135168 -6912 135494 -6910
rect 137704 -6912 138540 -6736
rect 135168 -8401 138540 -6912
rect 138356 -8719 138546 -8689
rect 138356 -9858 138379 -8719
rect 138540 -9858 138546 -8719
rect 138356 -9889 138546 -9858
use bias_nstack  bias_nstack_0
array 0 75 -534 0 0 -4355
timestamp 1717035242
transform 1 0 133578 0 -1 18020
box 3258 -2860 3926 1035
use bias_nstack  bias_nstack_1
array 0 87 -534 0 0 -4355
timestamp 1717035242
transform -1 0 94395 0 -1 8820
box 3258 -2860 3926 1035
use bias_nstack  bias_nstack_2
array 0 87 -534 0 0 -4355
timestamp 1717035242
transform -1 0 94395 0 -1 -380
box 3258 -2860 3926 1035
use bias_nstack  bias_nstack_3
array 0 3 -534 0 0 -4355
timestamp 1717035242
transform -1 0 139251 0 -1 -9580
box 3258 -2860 3926 1035
use bias_pstack  bias_pstack_0
array 0 75 534 0 0 -4355
timestamp 1717035242
transform -1 0 139531 0 -1 21426
box 1986 -3967 2714 388
use bias_pstack  bias_pstack_1
array 0 87 534 0 0 -4355
timestamp 1717035242
transform 1 0 88442 0 -1 12226
box 1986 -3967 2714 388
use bias_pstack  bias_pstack_2
array 0 87 534 0 0 -4355
timestamp 1717035242
transform 1 0 88442 0 -1 3026
box 1986 -3967 2714 388
use bias_pstack  bias_pstack_3
array 0 3 534 0 0 -4355
timestamp 1717035242
transform 1 0 133298 0 -1 -6174
box 1986 -3967 2714 388
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_8 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform 1 0 91893 0 1 17858
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_9
timestamp 1715205430
transform 1 0 91893 0 1 21114
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_10
timestamp 1715205430
transform 1 0 91893 0 1 19486
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_11
timestamp 1715205430
transform 1 0 94485 0 1 17858
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_12
timestamp 1715205430
transform 1 0 91893 0 1 22742
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_13
timestamp 1715205430
transform 1 0 94485 0 1 22742
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_16
timestamp 1715205430
transform 1 0 94485 0 1 21114
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_17
timestamp 1715205430
transform 1 0 94485 0 1 19486
box -66 -43 450 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_8 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform 1 0 92277 0 1 17858
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_9
timestamp 1715205430
transform 1 0 92277 0 1 21114
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_10
timestamp 1715205430
transform 1 0 92277 0 1 19486
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_11
timestamp 1715205430
transform 1 0 94869 0 1 17858
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_12
timestamp 1715205430
transform 1 0 92277 0 1 22742
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_13
timestamp 1715205430
transform 1 0 94869 0 1 22742
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_16
timestamp 1715205430
transform 1 0 94869 0 1 21114
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_17
timestamp 1715205430
transform 1 0 94869 0 1 19486
box -66 -43 162 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform 1 0 94485 0 -1 19486
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_1
timestamp 1715205430
transform 1 0 91893 0 -1 19486
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_2
timestamp 1715205430
transform 1 0 94485 0 -1 21114
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_3
timestamp 1715205430
transform 1 0 94485 0 -1 22742
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_4
timestamp 1715205430
transform 1 0 91893 0 -1 24370
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_7
timestamp 1715205430
transform 1 0 91893 0 -1 21114
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_10
timestamp 1715205430
transform 1 0 94485 0 -1 24370
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_11
timestamp 1715205430
transform 1 0 91893 0 -1 22742
box -66 -43 546 897
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
array 0 1 -2592 0 3 1628
timestamp 1715205430
transform 1 0 92373 0 1 17858
box -66 -43 2178 1671
<< labels >>
flabel metal4 135168 -8401 135401 -6716 0 FreeSans 1600 90 0 0 avss
port 2 nsew
flabel metal4 135167 -6565 135400 -4880 0 FreeSans 1600 90 0 0 avdd
port 1 nsew
flabel metal4 90311 2635 90544 4320 0 FreeSans 1600 90 0 0 avdd
port 1 nsew
flabel metal4 90312 799 90545 2484 0 FreeSans 1600 90 0 0 avss
port 2 nsew
flabel metal4 90311 11835 90544 13520 0 FreeSans 1600 90 0 0 avdd
port 1 nsew
flabel metal4 90312 9999 90545 11684 0 FreeSans 1600 90 0 0 avss
port 2 nsew
flabel metal4 137603 21035 137662 22720 0 FreeSans 1600 90 0 0 avdd
port 1 nsew
flabel metal4 137603 19199 137661 20884 0 FreeSans 1600 90 0 0 avss
port 2 nsew
flabel metal4 88136 23083 88736 24283 0 FreeSans 3200 90 0 0 dvdd
port 3 nsew
flabel metal4 88136 21035 88736 22720 0 FreeSans 3200 90 0 0 avdd
port 1 nsew
flabel metal4 88136 19199 88736 20884 0 FreeSans 3200 90 0 0 avss
port 2 nsew
flabel metal4 88136 17711 88736 18911 0 FreeSans 3200 90 0 0 dvss
port 4 nsew
flabel metal2 92702 17078 92742 17478 0 FreeSans 400 90 0 0 en_snk_test
port 26 nsew
flabel metal2 92578 17078 92618 17453 0 FreeSans 400 90 0 0 en_user2_trim_n
port 16 nsew
flabel metal2 92462 17078 92502 17453 0 FreeSans 400 90 0 0 en_comp_trim_n
port 24 nsew
flabel metal2 92342 17078 92382 17453 0 FreeSans 400 90 0 0 en_hsxo_trim_n
port 25 nsew
flabel metal2 90110 17078 90150 17453 0 FreeSans 400 90 0 0 en_lp2_bias
port 20 nsew
flabel metal2 89990 17078 90030 17453 0 FreeSans 400 90 0 0 en_lp1_trim_p
port 21 nsew
flabel metal2 89870 17078 89910 17453 0 FreeSans 400 90 0 0 en_lsxo_bias
port 23 nsew
flabel metal2 89750 17078 89790 17453 0 FreeSans 400 90 0 0 en_lp1_bias
port 22 nsew
<< end >>
