magic
tech sky130A
magscale 1 2
timestamp 1716925370
<< error_p >>
rect 20242 6143 20244 7195
rect 20036 5937 20450 6143
rect 20036 5935 21502 5937
rect 20036 5729 20450 5935
<< error_s >>
rect 44269 8352 47212 8386
rect 41597 8142 49898 8176
rect 41597 4236 49898 4409
rect 41597 3870 49898 4043
rect 41597 278 49898 312
rect 41597 46 49898 105
use bias_generator_be  bias_generator_be_0
timestamp 1716920177
transform 1 0 45529 0 1 -418
box 0 0 152006 9467
use bias_generator_fe  bias_generator_fe_0
timestamp 1716925370
transform 1 0 0 0 1 0
box 1072 0 45966 8863
<< end >>
