magic
tech sky130A
magscale 1 2
timestamp 1717106147
<< error_s >>
rect -24 925 876 1825
<< dnwell >>
rect -24 719 138229 8571
<< nwell >>
rect -24 8365 138338 8680
rect 138023 925 138338 8365
rect -24 610 138338 925
<< pwell >>
rect 2095 925 2183 947
<< mvpsubdiff >>
rect 42 8770 327 8804
rect 138398 8770 138458 8804
rect 138424 8744 138458 8770
rect 139072 8182 139132 8216
rect 149416 8182 149476 8216
rect 139072 8156 139106 8182
rect 139072 1252 139106 1278
rect 149442 8156 149476 8182
rect 149442 1252 149476 1278
rect 139072 1218 139132 1252
rect 149416 1218 149476 1252
rect 138424 498 138458 524
rect 42 464 299 498
rect 138398 464 138458 498
<< mvnsubdiff >>
rect 42 8594 138272 8614
rect 42 8560 327 8594
rect 138192 8560 138272 8594
rect 42 8540 138272 8560
rect 138198 8534 138272 8540
rect 138198 756 138218 8534
rect 138252 756 138272 8534
rect 138198 750 138272 756
rect 42 730 138272 750
rect 42 696 299 730
rect 138192 696 138272 730
rect 42 676 138272 696
<< mvpsubdiffcont >>
rect 327 8770 138398 8804
rect 138424 524 138458 8744
rect 139132 8182 149416 8216
rect 139072 1278 139106 8156
rect 149442 1278 149476 8156
rect 139132 1218 149416 1252
rect 299 464 138398 498
<< mvnsubdiffcont >>
rect 327 8560 138192 8594
rect 138218 756 138252 8534
rect 299 696 138192 730
<< locali >>
rect 42 8770 327 8804
rect 138398 8770 138458 8804
rect 42 8755 138458 8770
rect 42 8671 138360 8755
rect 50 8560 327 8594
rect 138192 8560 138252 8594
rect 50 8534 138252 8560
rect 50 8529 138218 8534
rect 50 8375 138128 8529
rect 138081 909 138128 8375
rect 42 752 138128 909
rect 138187 756 138218 8529
rect 138187 752 138252 756
rect 42 730 138252 752
rect 42 696 299 730
rect 138192 696 138252 730
rect 138316 610 138360 8671
rect 42 523 138360 610
rect 42 464 299 523
rect 138307 514 138360 523
rect 138412 8744 138458 8755
rect 138412 524 138424 8744
rect 138458 8182 139132 8216
rect 149416 8182 149476 8216
rect 138458 8156 149476 8182
rect 138458 8019 139072 8156
rect 138458 1278 139072 1414
rect 139106 8094 149442 8156
rect 139106 1340 139189 8094
rect 141863 7594 141910 7660
rect 144455 7594 144502 7660
rect 147047 7594 147094 7660
rect 140909 6766 141079 6782
rect 140909 6664 140925 6766
rect 141058 6664 141079 6766
rect 140909 6648 141079 6664
rect 143501 6766 143671 6782
rect 143501 6664 143517 6766
rect 143650 6664 143671 6766
rect 143501 6648 143671 6664
rect 146093 6766 146263 6782
rect 146093 6664 146109 6766
rect 146242 6664 146263 6766
rect 146093 6648 146263 6664
rect 148685 6766 148855 6782
rect 148685 6664 148701 6766
rect 148834 6664 148855 6766
rect 148685 6648 148855 6664
rect 141863 5966 141910 6032
rect 144455 5966 144502 6032
rect 147047 5966 147094 6032
rect 140909 5138 141079 5154
rect 140909 5036 140925 5138
rect 141058 5036 141079 5138
rect 140909 5020 141079 5036
rect 143501 5138 143671 5154
rect 143501 5036 143517 5138
rect 143650 5036 143671 5138
rect 143501 5020 143671 5036
rect 146093 5138 146263 5154
rect 146093 5036 146109 5138
rect 146242 5036 146263 5138
rect 146093 5020 146263 5036
rect 148685 5138 148855 5154
rect 148685 5036 148701 5138
rect 148834 5036 148855 5138
rect 148685 5020 148855 5036
rect 144455 4338 144502 4404
rect 147047 4338 147094 4404
rect 140909 3510 141079 3526
rect 140909 3408 140925 3510
rect 141058 3408 141079 3510
rect 140909 3392 141079 3408
rect 143501 3510 143671 3526
rect 143501 3408 143517 3510
rect 143650 3408 143671 3510
rect 143501 3392 143671 3408
rect 146093 3510 146263 3526
rect 146093 3408 146109 3510
rect 146242 3408 146263 3510
rect 146093 3392 146263 3408
rect 148685 3510 148855 3526
rect 148685 3408 148701 3510
rect 148834 3408 148855 3510
rect 148685 3392 148855 3408
rect 144455 2710 144502 2776
rect 147047 2710 147094 2776
rect 140909 1882 141079 1898
rect 140909 1780 140925 1882
rect 141058 1780 141079 1882
rect 140909 1764 141079 1780
rect 143501 1882 143671 1898
rect 143501 1780 143517 1882
rect 143650 1780 143671 1882
rect 143501 1764 143671 1780
rect 146093 1882 146263 1898
rect 146093 1780 146109 1882
rect 146242 1780 146263 1882
rect 146093 1764 146263 1780
rect 148685 1882 148855 1898
rect 148685 1780 148701 1882
rect 148834 1780 148855 1882
rect 148685 1764 148855 1780
rect 149348 1340 149442 8094
rect 139106 1278 149442 1340
rect 138458 1252 149476 1278
rect 138458 1218 139132 1252
rect 149416 1218 149476 1252
rect 138458 1217 139161 1218
rect 138412 514 138458 524
rect 138307 498 138458 514
rect 138398 464 138458 498
<< viali >>
rect 138128 752 138187 8529
rect 299 498 138307 523
rect 138360 514 138412 8755
rect 141529 7624 141575 7803
rect 144121 7624 144167 7803
rect 146713 7624 146759 7803
rect 139318 7316 139366 7547
rect 140925 6664 141058 6766
rect 143517 6664 143650 6766
rect 146109 6664 146242 6766
rect 148701 6664 148834 6766
rect 141529 5996 141575 6175
rect 144121 5996 144167 6175
rect 146713 5996 146759 6175
rect 139318 5688 139366 5919
rect 140925 5036 141058 5138
rect 143517 5036 143650 5138
rect 146109 5036 146242 5138
rect 148701 5036 148834 5138
rect 144121 4368 144167 4547
rect 146713 4368 146759 4547
rect 139318 4060 139366 4291
rect 141910 4060 141958 4291
rect 140925 3408 141058 3510
rect 143517 3408 143650 3510
rect 146109 3408 146242 3510
rect 148701 3408 148834 3510
rect 144121 2740 144167 2919
rect 146713 2740 146759 2919
rect 139318 2432 139366 2663
rect 141910 2432 141958 2663
rect 140925 1780 141058 1882
rect 143517 1780 143650 1882
rect 146109 1780 146242 1882
rect 148701 1780 148834 1882
rect 299 479 138307 498
<< metal1 >>
rect 138332 8755 138448 8797
rect 138093 8529 138231 8580
rect 138093 6299 138128 8529
rect 138187 6299 138231 8529
rect 138093 4657 138108 6299
rect 138215 4657 138231 6299
rect 138093 752 138128 4657
rect 138187 752 138231 4657
rect 138093 705 138231 752
rect 138332 542 138360 8755
rect 138412 2512 138448 8755
rect 139317 8031 149260 8045
rect 139317 7872 142015 8031
rect 143290 7872 149260 8031
rect 141512 7815 141576 7816
rect 144108 7815 144172 7816
rect 141512 7814 141581 7815
rect 141512 7784 141518 7814
rect 141570 7803 141581 7814
rect 141472 7744 141518 7784
rect 141512 7614 141518 7744
rect 141575 7624 141581 7803
rect 141570 7614 141581 7624
rect 144108 7814 144173 7815
rect 144108 7614 144114 7814
rect 144166 7803 144173 7814
rect 144167 7624 144173 7803
rect 144166 7614 144173 7624
rect 141522 7612 141581 7614
rect 144114 7612 144173 7614
rect 146704 7814 146768 7816
rect 146704 7614 146710 7814
rect 146762 7614 146768 7814
rect 146704 7612 146768 7614
rect 139306 7547 139384 7553
rect 139306 7544 139318 7547
rect 139288 7542 139318 7544
rect 139288 7504 139314 7542
rect 139306 7342 139314 7504
rect 139306 7316 139318 7342
rect 139366 7316 139384 7547
rect 144132 7529 144172 7612
rect 146720 7600 146760 7612
rect 139306 7310 139384 7316
rect 139306 7066 144593 7239
rect 145872 7066 149249 7239
rect 141028 6946 147328 7003
rect 140909 6766 141079 6782
rect 140909 6664 140925 6766
rect 141058 6664 141079 6766
rect 140909 6648 141079 6664
rect 143501 6766 143671 6782
rect 143501 6664 143517 6766
rect 143650 6664 143671 6766
rect 143501 6648 143671 6664
rect 146093 6766 146263 6782
rect 146093 6664 146109 6766
rect 146242 6664 146263 6766
rect 146093 6648 146263 6664
rect 148685 6766 148855 6782
rect 148685 6664 148701 6766
rect 148834 6664 148855 6766
rect 148685 6648 148855 6664
rect 139306 6249 142018 6422
rect 143288 6249 149249 6422
rect 141512 6187 141576 6188
rect 141512 6186 141581 6187
rect 141512 6156 141518 6186
rect 141570 6175 141581 6186
rect 141482 6116 141518 6156
rect 141512 5986 141518 6116
rect 141575 5996 141581 6175
rect 141570 5986 141581 5996
rect 144108 6186 144174 6188
rect 146706 6186 146765 6187
rect 144108 5986 144114 6186
rect 144166 6175 144174 6186
rect 144167 5996 144174 6175
rect 144166 5986 144174 5996
rect 146704 5986 146710 6186
rect 146762 5986 146768 6186
rect 141522 5984 141581 5986
rect 144114 5984 144173 5986
rect 146704 5984 146768 5986
rect 139306 5919 139384 5925
rect 139306 5916 139318 5919
rect 139288 5914 139318 5916
rect 139288 5876 139314 5914
rect 139306 5714 139314 5876
rect 139306 5688 139318 5714
rect 139366 5688 139384 5919
rect 144132 5901 144172 5984
rect 146720 5980 146760 5984
rect 139306 5682 139384 5688
rect 139323 5438 144589 5611
rect 145868 5438 149266 5611
rect 140862 5318 147328 5375
rect 140909 5138 141079 5154
rect 140909 5036 140925 5138
rect 141058 5036 141079 5138
rect 140909 5020 141079 5036
rect 143501 5138 143671 5154
rect 143501 5036 143517 5138
rect 143650 5036 143671 5138
rect 143501 5020 143671 5036
rect 146093 5138 146263 5154
rect 146093 5036 146109 5138
rect 146242 5036 146263 5138
rect 146093 5020 146263 5036
rect 148685 5138 148855 5154
rect 148685 5036 148701 5138
rect 148834 5036 148855 5138
rect 148685 5020 148855 5036
rect 139295 4622 142016 4795
rect 143286 4622 149238 4795
rect 144108 4559 144172 4560
rect 144108 4558 144173 4559
rect 146706 4558 146765 4559
rect 144108 4528 144114 4558
rect 144166 4547 144173 4558
rect 138822 4168 138828 4368
rect 138880 4328 141959 4368
rect 144108 4358 144114 4488
rect 144167 4368 144173 4547
rect 144166 4358 144173 4368
rect 144114 4356 144173 4358
rect 146704 4358 146710 4558
rect 146762 4358 146768 4558
rect 146704 4356 146768 4358
rect 146720 4350 146760 4356
rect 138880 4168 138886 4328
rect 141919 4297 141959 4328
rect 139306 4291 139384 4297
rect 139306 4288 139318 4291
rect 139288 4286 139318 4288
rect 139288 4248 139314 4286
rect 139306 4086 139314 4248
rect 139306 4060 139318 4086
rect 139366 4060 139384 4291
rect 139306 4054 139384 4060
rect 141898 4291 141974 4297
rect 141898 4060 141910 4291
rect 141958 4060 141974 4291
rect 141898 4054 141974 4060
rect 139312 3822 144593 3995
rect 145872 3822 149255 3995
rect 140689 3690 147328 3747
rect 140909 3510 141079 3526
rect 140909 3408 140925 3510
rect 141058 3408 141079 3510
rect 140909 3392 141079 3408
rect 143501 3510 143671 3526
rect 143501 3408 143517 3510
rect 143650 3408 143671 3510
rect 143501 3392 143671 3408
rect 146093 3510 146263 3526
rect 146093 3408 146109 3510
rect 146242 3408 146263 3510
rect 146093 3392 146263 3408
rect 148685 3510 148855 3526
rect 148685 3408 148701 3510
rect 148834 3408 148855 3510
rect 148685 3392 148855 3408
rect 139279 3000 142020 3173
rect 143290 3000 149222 3173
rect 144108 2930 144174 2932
rect 146706 2930 146765 2931
rect 144108 2900 144114 2930
rect 144166 2919 144174 2930
rect 138932 2540 138938 2740
rect 138990 2700 141955 2740
rect 144108 2730 144114 2860
rect 144167 2740 144174 2919
rect 144166 2730 144174 2740
rect 146704 2730 146710 2930
rect 146762 2730 146768 2930
rect 144114 2728 144173 2730
rect 146704 2728 146768 2730
rect 146720 2710 146760 2728
rect 138990 2540 138996 2700
rect 141915 2669 141955 2700
rect 139306 2663 139384 2669
rect 139306 2660 139318 2663
rect 139288 2658 139318 2660
rect 139288 2620 139314 2658
rect 138412 2481 138622 2512
rect 138593 1342 138622 2481
rect 139306 2458 139314 2620
rect 139306 2432 139318 2458
rect 139366 2432 139384 2663
rect 139306 2426 139384 2432
rect 141898 2663 141971 2669
rect 141898 2432 141910 2663
rect 141958 2432 141971 2663
rect 141898 2426 141971 2432
rect 139323 2183 144593 2356
rect 145872 2183 149266 2356
rect 140862 2062 147328 2119
rect 140909 1882 141079 1898
rect 140909 1780 140925 1882
rect 141058 1780 141079 1882
rect 140909 1764 141079 1780
rect 143501 1882 143671 1898
rect 143501 1780 143517 1882
rect 143650 1780 143671 1882
rect 143501 1764 143671 1780
rect 146093 1882 146263 1898
rect 146093 1780 146109 1882
rect 146242 1780 146263 1882
rect 146093 1764 146263 1780
rect 148685 1882 148855 1898
rect 148685 1780 148701 1882
rect 148834 1780 148855 1882
rect 148685 1764 148855 1780
rect 139301 1461 142013 1539
rect 143285 1461 149188 1539
rect 42 523 138360 542
rect 42 479 299 523
rect 138307 514 138360 523
rect 138412 1310 138622 1342
rect 138412 514 138448 1310
rect 138307 479 138448 514
rect 42 464 138448 479
<< via1 >>
rect 138108 4657 138128 6299
rect 138128 4657 138187 6299
rect 138187 4657 138215 6299
rect 142015 7868 143290 8031
rect 141518 7803 141570 7814
rect 141518 7624 141529 7803
rect 141529 7624 141570 7803
rect 141518 7614 141570 7624
rect 144114 7803 144166 7814
rect 144114 7624 144121 7803
rect 144121 7624 144166 7803
rect 144114 7614 144166 7624
rect 146710 7803 146762 7814
rect 146710 7624 146713 7803
rect 146713 7624 146759 7803
rect 146759 7624 146762 7803
rect 146710 7614 146762 7624
rect 139314 7342 139318 7542
rect 139318 7342 139366 7542
rect 144593 7047 145872 7264
rect 147328 6946 148322 7003
rect 140925 6664 141058 6766
rect 143517 6664 143650 6766
rect 146109 6664 146242 6766
rect 148701 6664 148834 6766
rect 142018 6229 143288 6444
rect 141518 6175 141570 6186
rect 141518 5996 141529 6175
rect 141529 5996 141570 6175
rect 141518 5986 141570 5996
rect 144114 6175 144166 6186
rect 144114 5996 144121 6175
rect 144121 5996 144166 6175
rect 144114 5986 144166 5996
rect 146710 6175 146762 6186
rect 146710 5996 146713 6175
rect 146713 5996 146759 6175
rect 146759 5996 146762 6175
rect 146710 5986 146762 5996
rect 139314 5714 139318 5914
rect 139318 5714 139366 5914
rect 144589 5420 145868 5637
rect 147328 5318 148322 5375
rect 140925 5036 141058 5138
rect 143517 5036 143650 5138
rect 146109 5036 146242 5138
rect 148701 5036 148834 5138
rect 142016 4609 143286 4824
rect 144114 4547 144166 4558
rect 138828 4168 138880 4368
rect 144114 4368 144121 4547
rect 144121 4368 144166 4547
rect 144114 4358 144166 4368
rect 146710 4547 146762 4558
rect 146710 4368 146713 4547
rect 146713 4368 146759 4547
rect 146759 4368 146762 4547
rect 146710 4358 146762 4368
rect 139314 4086 139318 4286
rect 139318 4086 139366 4286
rect 144593 3789 145872 4006
rect 147328 3690 148322 3747
rect 140925 3408 141058 3510
rect 143517 3408 143650 3510
rect 146109 3408 146242 3510
rect 148701 3408 148834 3510
rect 142020 2976 143290 3191
rect 144114 2919 144166 2930
rect 138938 2540 138990 2740
rect 144114 2740 144121 2919
rect 144121 2740 144166 2919
rect 144114 2730 144166 2740
rect 146710 2919 146762 2930
rect 146710 2740 146713 2919
rect 146713 2740 146759 2919
rect 146759 2740 146762 2919
rect 146710 2730 146762 2740
rect 138379 1342 138412 2481
rect 138412 1342 138593 2481
rect 139314 2458 139318 2658
rect 139318 2458 139366 2658
rect 144593 2163 145872 2380
rect 147328 2062 148322 2119
rect 140925 1780 141058 1882
rect 143517 1780 143650 1882
rect 146109 1780 146242 1882
rect 148701 1780 148834 1882
rect 142013 1448 143285 1563
<< metal2 >>
rect 127394 9730 147076 9778
rect 127394 9346 127442 9730
rect 117318 9298 127442 9346
rect 127550 9634 146890 9682
rect 117318 9138 117366 9298
rect 127550 9254 127598 9634
rect 106814 9090 117366 9138
rect 117506 9206 127598 9254
rect 127696 9538 146756 9586
rect 33557 8967 33725 8969
rect 331 8737 41568 8967
rect 331 8735 33557 8737
rect 33725 8735 41568 8737
rect 41887 8735 106714 8967
rect 106814 8660 106862 9090
rect 107110 8735 112834 8967
rect 113161 8735 117368 8967
rect 117506 8660 117554 9206
rect 127696 9134 127744 9538
rect 123920 9086 127744 9134
rect 128202 9442 146620 9490
rect 117754 8735 121402 8967
rect 121729 8735 123820 8967
rect 123920 8660 123968 9086
rect 124170 8735 126662 8967
rect 126989 8735 128064 8967
rect 128202 8660 128250 9442
rect 130336 9346 144478 9394
rect 128539 8735 129832 8967
rect 130159 8735 130186 8967
rect 130336 8660 130384 9346
rect 134516 9250 144322 9298
rect 134516 9114 134564 9250
rect 132658 9066 134564 9114
rect 134708 9154 144160 9202
rect 130685 8735 131924 8967
rect 132251 8735 132590 8967
rect 132658 8660 132706 9066
rect 132825 8735 134016 8967
rect 134343 8735 134640 8967
rect 134708 8660 134756 9154
rect 517 8428 40683 8660
rect 40866 8428 106872 8660
rect 107270 8428 111939 8660
rect 112124 8428 117562 8660
rect 117926 8428 120507 8660
rect 120692 8428 123968 8660
rect 124197 8428 125767 8660
rect 125952 8428 128250 8660
rect 128617 8428 128937 8660
rect 129122 8428 130384 8660
rect 130721 8428 131029 8660
rect 131214 8612 132706 8660
rect 131214 8428 132590 8612
rect 132825 8428 133121 8660
rect 133306 8612 134756 8660
rect 134812 9058 144012 9106
rect 134812 8658 134860 9058
rect 134929 8735 135568 8967
rect 135895 8735 135909 8967
rect 135981 8735 135997 8967
rect 136169 8735 136203 8967
rect 136506 8735 136678 8967
rect 136895 8735 137113 8967
rect 134929 8658 135213 8660
rect 133306 8428 134640 8612
rect 134812 8610 135213 8658
rect 134929 8428 135213 8610
rect 135398 8428 135858 8660
rect 135981 8428 136339 8660
rect 136524 8428 136549 8660
rect 136693 8428 137022 8660
rect 137197 8520 137292 8660
rect 137197 8480 141564 8520
rect 137197 8428 137292 8480
rect 136494 8372 136534 8428
rect 141354 8372 141394 8376
rect 136494 8332 141394 8372
rect 66 8027 137616 8265
rect 66 7696 188 7930
rect 137608 7696 137655 7930
rect 137910 7696 137939 7930
rect 139320 7552 139360 8012
rect 139314 7542 139366 7552
rect 141354 7384 141394 8332
rect 141524 7824 141564 8480
rect 142000 8031 143303 8086
rect 142000 7868 142015 8031
rect 143290 7868 143303 8031
rect 141518 7814 141570 7824
rect 141518 7606 141570 7614
rect 141354 7344 141564 7384
rect 139314 7334 139366 7342
rect 139320 6982 139360 7334
rect 139320 6942 139748 6982
rect 66 6696 137616 6930
rect 66 6695 186 6696
rect 138079 6299 138270 6322
rect 182 5692 137616 5926
rect 317 4654 392 4738
rect 137608 4638 137654 4872
rect 137909 4638 137938 4872
rect 138079 4657 138108 6299
rect 138215 4657 138270 6299
rect 139320 5924 139360 6384
rect 139314 5914 139366 5924
rect 139314 5706 139366 5714
rect 139320 4904 139360 5706
rect 139320 4864 139616 4904
rect 138079 4638 138270 4657
rect 66 4461 1279 4480
rect 66 4377 392 4461
rect 66 4242 1279 4377
rect 138828 4368 138880 4376
rect 139320 4296 139360 4756
rect 138828 4162 138880 4168
rect 139314 4286 139366 4296
rect 223 3218 137597 3456
rect 138358 2481 138622 2512
rect 165 2234 137589 2472
rect 66 1246 137597 1484
rect 138358 1342 138379 2481
rect 138593 1342 138622 2481
rect 138358 1310 138622 1342
rect 138834 1172 138874 4162
rect 139314 4078 139366 4086
rect 139320 3294 139360 4078
rect 139320 3254 139488 3294
rect 138938 2740 138990 2748
rect 139320 2668 139360 3128
rect 138938 2534 138990 2540
rect 139314 2658 139366 2668
rect 136210 1132 138874 1172
rect 136210 1037 136250 1132
rect 66 849 36216 1037
rect 36401 849 74838 1037
rect 75258 1020 96188 1037
rect 75258 858 85718 1020
rect 85914 858 96188 1020
rect 75258 849 96188 858
rect 96610 849 105496 1037
rect 105681 849 117562 1037
rect 117942 849 120004 1037
rect 120189 849 128242 1037
rect 128654 849 135068 1037
rect 135185 849 136250 1037
rect 136690 849 137068 1037
rect 137185 972 137300 1037
rect 138944 972 138984 2534
rect 139314 2450 139366 2458
rect 137185 932 138984 972
rect 137185 849 137300 932
rect 66 593 37111 781
rect 37438 593 74676 781
rect 74776 342 74824 849
rect 75096 768 96022 781
rect 75096 608 86620 768
rect 86946 608 96022 768
rect 75096 593 96022 608
rect 96130 466 96178 849
rect 96444 593 106391 781
rect 106718 593 117400 781
rect 96130 418 117026 466
rect 74776 294 116876 342
rect 116978 326 117026 418
rect 117496 422 117544 849
rect 117780 593 120899 781
rect 121226 593 128070 781
rect 128194 518 128242 849
rect 128482 593 134680 781
rect 134862 593 136081 781
rect 136525 593 136680 781
rect 136862 593 137135 781
rect 139320 518 139360 2450
rect 128194 470 139360 518
rect 139448 422 139488 3254
rect 117496 374 139488 422
rect 139576 326 139616 4864
rect 116828 230 116876 294
rect 116972 278 139616 326
rect 139708 230 139748 6942
rect 140909 6766 141079 6782
rect 140909 6664 140925 6766
rect 141058 6739 141079 6766
rect 141058 6699 141439 6739
rect 141058 6664 141079 6699
rect 140909 6648 141079 6664
rect 140909 5138 141079 5154
rect 140909 5036 140925 5138
rect 141058 5097 141079 5138
rect 141058 5057 141319 5097
rect 141058 5036 141079 5057
rect 140909 5020 141079 5036
rect 140909 3510 141079 3526
rect 140909 3408 140925 3510
rect 141058 3474 141079 3510
rect 141058 3434 141199 3474
rect 141058 3408 141079 3434
rect 140909 3392 141079 3408
rect 140909 1882 141079 1898
rect 140909 1780 140925 1882
rect 141058 1780 141079 1882
rect 140909 1764 141079 1780
rect 141039 678 141079 1764
rect 141159 678 141199 3434
rect 141279 678 141319 5057
rect 141399 678 141439 6699
rect 141524 6196 141564 7344
rect 142000 6444 143303 7868
rect 143972 7194 144012 9058
rect 144120 7824 144160 9154
rect 144114 7814 144166 7824
rect 144114 7606 144166 7614
rect 143972 7154 144160 7194
rect 143501 6766 143671 6782
rect 143501 6664 143517 6766
rect 143650 6739 143671 6766
rect 143650 6699 144031 6739
rect 143650 6664 143671 6699
rect 143501 6648 143671 6664
rect 142000 6229 142018 6444
rect 143288 6229 143303 6444
rect 141518 6186 141570 6196
rect 141518 5978 141570 5986
rect 142000 4824 143303 6229
rect 143501 5138 143671 5154
rect 143501 5036 143517 5138
rect 143650 5097 143671 5138
rect 143650 5057 143911 5097
rect 143650 5036 143671 5057
rect 143501 5020 143671 5036
rect 142000 4609 142016 4824
rect 143286 4609 143303 4824
rect 142000 3191 143303 4609
rect 143501 3510 143671 3526
rect 143501 3408 143517 3510
rect 143650 3474 143671 3510
rect 143650 3434 143791 3474
rect 143650 3408 143671 3434
rect 143501 3392 143671 3408
rect 142000 2976 142020 3191
rect 143290 2976 143303 3191
rect 142000 2485 143303 2976
rect 142000 1563 142027 2485
rect 143269 1563 143303 2485
rect 143501 1882 143671 1898
rect 143501 1780 143517 1882
rect 143650 1780 143671 1882
rect 143501 1764 143671 1780
rect 142000 1448 142013 1563
rect 143285 1448 143303 1563
rect 142000 1340 142027 1448
rect 143269 1340 143303 1448
rect 142000 1300 143303 1340
rect 143631 678 143671 1764
rect 143751 678 143791 3434
rect 143871 678 143911 5057
rect 143991 678 144031 6699
rect 144120 6196 144160 7154
rect 144114 6186 144166 6196
rect 144114 5978 144166 5986
rect 144282 5302 144322 9250
rect 144120 5262 144322 5302
rect 144120 4568 144160 5262
rect 144114 4558 144166 4568
rect 144114 4350 144166 4358
rect 144438 4076 144478 9346
rect 144120 4036 144478 4076
rect 144580 7264 145885 8101
rect 144580 7047 144593 7264
rect 145872 7047 145885 7264
rect 146580 7178 146620 9442
rect 146716 7824 146756 9538
rect 146710 7814 146762 7824
rect 146710 7606 146762 7614
rect 146580 7138 146756 7178
rect 144580 6280 145885 7047
rect 146093 6766 146263 6782
rect 146093 6664 146109 6766
rect 146242 6739 146263 6766
rect 146242 6699 146623 6739
rect 146242 6664 146263 6699
rect 146093 6648 146263 6664
rect 144580 5637 144639 6280
rect 145841 5637 145885 6280
rect 144580 5420 144589 5637
rect 145868 5420 145885 5637
rect 144580 4689 144639 5420
rect 145841 4689 145885 5420
rect 146093 5138 146263 5154
rect 146093 5036 146109 5138
rect 146242 5097 146263 5138
rect 146242 5057 146503 5097
rect 146242 5036 146263 5057
rect 146093 5020 146263 5036
rect 144120 2940 144160 4036
rect 144580 4006 145885 4689
rect 144580 3789 144593 4006
rect 145872 3789 145885 4006
rect 144114 2930 144166 2940
rect 144114 2722 144166 2730
rect 144580 2380 145885 3789
rect 146093 3510 146263 3526
rect 146093 3408 146109 3510
rect 146242 3474 146263 3510
rect 146242 3434 146383 3474
rect 146242 3408 146263 3434
rect 146093 3392 146263 3408
rect 144580 2163 144593 2380
rect 145872 2163 145885 2380
rect 144580 1390 145885 2163
rect 146093 1882 146263 1898
rect 146093 1780 146109 1882
rect 146242 1780 146263 1882
rect 146093 1764 146263 1780
rect 146223 678 146263 1764
rect 146343 678 146383 3434
rect 146463 678 146503 5057
rect 146583 678 146623 6699
rect 146716 6196 146756 7138
rect 146710 6186 146762 6196
rect 146710 5978 146762 5986
rect 146850 5870 146890 9634
rect 146716 5830 146890 5870
rect 146716 4568 146756 5830
rect 146710 4558 146762 4568
rect 146710 4350 146762 4358
rect 147036 4090 147076 9730
rect 146716 4050 147076 4090
rect 147328 7851 148322 8094
rect 147328 7003 147359 7851
rect 148291 7003 148322 7851
rect 147328 6713 147359 6946
rect 148291 6713 148322 6946
rect 147328 5375 148322 6713
rect 148685 6766 148855 6782
rect 148685 6664 148701 6766
rect 148834 6739 148855 6766
rect 148834 6699 149215 6739
rect 148834 6664 148855 6699
rect 148685 6648 148855 6664
rect 146716 2940 146756 4050
rect 147328 3747 148322 5318
rect 148685 5138 148855 5154
rect 148685 5036 148701 5138
rect 148834 5097 148855 5138
rect 148834 5057 149095 5097
rect 148834 5036 148855 5057
rect 148685 5020 148855 5036
rect 146710 2930 146762 2940
rect 146710 2722 146762 2730
rect 147328 2119 148322 3690
rect 148685 3510 148855 3526
rect 148685 3408 148701 3510
rect 148834 3474 148855 3510
rect 148834 3434 148975 3474
rect 148834 3408 148855 3434
rect 148685 3392 148855 3408
rect 147328 1301 148322 2062
rect 148685 1882 148855 1898
rect 148685 1780 148701 1882
rect 148834 1780 148855 1882
rect 148685 1764 148855 1780
rect 148815 678 148855 1764
rect 148935 678 148975 3434
rect 149055 678 149095 5057
rect 149175 678 149215 6699
rect 116828 182 139748 230
<< via2 >>
rect 41568 8735 41887 8967
rect 112834 8735 113161 8967
rect 121402 8735 121729 8967
rect 126662 8735 126989 8967
rect 129832 8735 130159 8967
rect 131924 8735 132251 8967
rect 134016 8735 134343 8967
rect 40683 8428 40866 8660
rect 111939 8428 112124 8660
rect 120507 8428 120692 8660
rect 125767 8428 125952 8660
rect 128937 8428 129122 8660
rect 131029 8428 131214 8660
rect 133121 8428 133306 8660
rect 135568 8735 135895 8967
rect 135997 8735 136169 8967
rect 136678 8735 136895 8967
rect 135213 8428 135398 8660
rect 136339 8428 136524 8660
rect 137022 8428 137197 8660
rect 137655 7696 137910 7930
rect 392 4654 33298 4738
rect 33715 4654 137146 4738
rect 137654 4638 137909 4872
rect 138108 4657 138215 6299
rect 392 4377 33299 4461
rect 33716 4379 137147 4463
rect 138379 1342 138593 2481
rect 36216 849 36401 1037
rect 85718 858 85914 1020
rect 105496 849 105681 1037
rect 120004 849 120189 1037
rect 135068 849 135185 1037
rect 137068 849 137185 1037
rect 37111 593 37438 781
rect 86620 608 86946 768
rect 106391 593 106718 781
rect 120899 593 121226 781
rect 134680 593 134862 781
rect 136680 593 136862 781
rect 142027 1563 143269 2485
rect 142027 1448 143269 1563
rect 142027 1340 143269 1448
rect 144639 5637 145841 6280
rect 144639 5420 145841 5637
rect 144639 4689 145841 5420
rect 147359 7003 148291 7851
rect 147359 6946 148291 7003
rect 147359 6713 148291 6946
<< metal3 >>
rect 40664 8660 40885 9465
rect 41542 8967 41905 9465
rect 41542 8735 41568 8967
rect 41887 8735 41905 8967
rect 41542 8714 41905 8735
rect 40664 8428 40683 8660
rect 40866 8428 40885 8660
rect 40664 8390 40885 8428
rect 111922 8660 112143 9465
rect 112817 8967 113179 9465
rect 112817 8735 112834 8967
rect 113161 8735 113179 8967
rect 112817 8714 113179 8735
rect 111922 8428 111939 8660
rect 112124 8428 112143 8660
rect 111922 8390 112143 8428
rect 120490 8660 120711 9466
rect 121385 8967 121747 9465
rect 121385 8735 121402 8967
rect 121729 8735 121747 8967
rect 121385 8714 121747 8735
rect 120490 8428 120507 8660
rect 120692 8428 120711 8660
rect 120490 8390 120711 8428
rect 125750 8660 125971 9465
rect 126645 8967 127003 9465
rect 126645 8735 126662 8967
rect 126989 8735 127003 8967
rect 126645 8714 127003 8735
rect 125750 8428 125767 8660
rect 125952 8428 125971 8660
rect 125750 8390 125971 8428
rect 128920 8660 129141 9465
rect 129815 8967 130173 9465
rect 129815 8735 129832 8967
rect 130159 8735 130173 8967
rect 129815 8714 130173 8735
rect 128920 8428 128937 8660
rect 129122 8428 129141 8660
rect 128920 8390 129141 8428
rect 131012 8660 131233 9465
rect 131907 8967 132265 9465
rect 131907 8735 131924 8967
rect 132251 8735 132265 8967
rect 131907 8714 132265 8735
rect 131012 8428 131029 8660
rect 131214 8428 131233 8660
rect 131012 8390 131233 8428
rect 133104 8660 133325 9465
rect 133999 8967 134357 9465
rect 133999 8735 134016 8967
rect 134343 8735 134357 8967
rect 133999 8714 134357 8735
rect 133104 8428 133121 8660
rect 133306 8428 133325 8660
rect 133104 8390 133325 8428
rect 135196 8660 135417 9465
rect 135551 8967 135909 9465
rect 135551 8735 135568 8967
rect 135895 8735 135909 8967
rect 135551 8714 135909 8735
rect 135980 8967 136219 9465
rect 135980 8735 135997 8967
rect 136169 8735 136219 8967
rect 135980 8714 136219 8735
rect 135196 8428 135213 8660
rect 135398 8428 135417 8660
rect 135196 8390 135417 8428
rect 136322 8660 136543 9465
rect 136664 8967 136907 9466
rect 136664 8735 136678 8967
rect 136895 8735 136907 8967
rect 136664 8715 136907 8735
rect 136322 8428 136339 8660
rect 136524 8428 136543 8660
rect 136322 8390 136543 8428
rect 137011 8660 137210 9467
rect 137011 8428 137022 8660
rect 137197 8428 137210 8660
rect 137011 8408 137210 8428
rect 137642 7930 137920 7967
rect 137642 7696 137655 7930
rect 137910 7696 137920 7930
rect 137642 4872 137920 7696
rect 147328 7851 148321 7886
rect 147328 6713 147359 7851
rect 148291 6713 148321 7851
rect 147328 6684 148321 6713
rect 292 4827 137654 4872
rect 292 4654 392 4827
rect 292 4653 33715 4654
rect 137147 4653 137654 4827
rect 292 4638 137654 4653
rect 137909 4638 137920 4872
rect 138079 6299 138248 6321
rect 138079 4657 138108 6299
rect 138215 4657 138248 6299
rect 138079 4638 138248 4657
rect 144580 6280 145886 6323
rect 144580 4689 144639 6280
rect 145841 4689 145886 6280
rect 279 4464 137539 4480
rect 279 4461 33715 4464
rect 279 4288 392 4461
rect 137147 4290 137539 4464
rect 33758 4288 137539 4290
rect 279 4242 137539 4288
rect 137642 1254 137920 4638
rect 144580 4636 145886 4689
rect 138358 2481 138622 2512
rect 138358 1342 138379 2481
rect 138593 1342 138622 2481
rect 138358 1310 138622 1342
rect 142001 2485 143301 2513
rect 142001 1340 142027 2485
rect 143269 1340 143301 2485
rect 142001 1313 143301 1340
rect 36199 1037 36420 1075
rect 36199 849 36216 1037
rect 36401 849 36420 1037
rect 36199 0 36420 849
rect 85706 1020 85927 1075
rect 85706 858 85718 1020
rect 85914 858 85927 1020
rect 37094 781 37456 802
rect 37094 593 37111 781
rect 37438 593 37456 781
rect 37094 0 37456 593
rect 85706 0 85927 858
rect 105479 1037 105700 1076
rect 105479 849 105496 1037
rect 105681 849 105700 1037
rect 86601 768 86963 802
rect 86601 608 86620 768
rect 86946 608 86963 768
rect 86601 0 86963 608
rect 105479 1 105700 849
rect 119987 1037 120208 1076
rect 119987 849 120004 1037
rect 120189 849 120208 1037
rect 106374 781 106736 803
rect 106374 593 106391 781
rect 106718 593 106736 781
rect 106374 1 106736 593
rect 119987 1 120208 849
rect 135060 1037 135194 1053
rect 135060 849 135068 1037
rect 135185 849 135194 1037
rect 120882 781 121244 803
rect 120882 593 120899 781
rect 121226 593 121244 781
rect 120882 1 121244 593
rect 134670 781 134875 800
rect 134670 593 134680 781
rect 134862 593 134875 781
rect 134670 193 134875 593
rect 135060 195 135194 849
rect 137060 1037 137194 1053
rect 137060 849 137068 1037
rect 137185 849 137194 1037
rect 136670 781 136875 800
rect 136670 593 136680 781
rect 136862 593 136875 781
rect 136670 193 136875 593
rect 137060 195 137194 849
<< via3 >>
rect 147359 6713 148291 7851
rect 392 4738 137147 4827
rect 392 4654 33298 4738
rect 33298 4654 33715 4738
rect 33715 4654 137146 4738
rect 137146 4654 137147 4738
rect 33715 4653 137147 4654
rect 138108 4657 138215 6299
rect 144639 4689 145841 6280
rect 33715 4463 137147 4464
rect 33715 4461 33716 4463
rect 392 4377 33299 4461
rect 33299 4379 33716 4461
rect 33716 4379 137147 4463
rect 33299 4377 137147 4379
rect 392 4290 137147 4377
rect 392 4288 33758 4290
rect 138379 1342 138593 2481
rect 142027 1340 143269 2485
<< metal4 >>
rect 138356 7851 149477 7883
rect 138356 6713 147359 7851
rect 148291 6713 149477 7851
rect 138356 6683 149477 6713
rect 65 6299 149477 6320
rect 65 4827 138108 6299
rect 65 4654 392 4827
rect 137147 4657 138108 4827
rect 138215 6280 149477 6299
rect 138215 4689 144639 6280
rect 145841 4689 149477 6280
rect 138215 4657 149477 4689
rect 65 4653 33715 4654
rect 137147 4653 149477 4657
rect 65 4635 149477 4653
rect 66 4464 149477 4484
rect 66 4461 33715 4464
rect 66 4288 392 4461
rect 137147 4290 149477 4464
rect 33758 4288 149477 4290
rect 66 2799 149477 4288
rect 138356 2485 149477 2511
rect 138356 2481 142027 2485
rect 138356 1342 138379 2481
rect 138593 1342 142027 2481
rect 138356 1340 142027 1342
rect 143269 1340 149477 2485
rect 138356 1311 149477 1340
use bias_nstack  bias_nstack_0
array 0 256 -534 0 0 -3895
timestamp 1717035242
transform -1 0 4149 0 -1 1620
box 3258 -2860 3926 1035
use bias_pstack  bias_pstack_0
array 0 256 534 0 0 -4355
timestamp 1717035242
transform 1 0 -1804 0 -1 5026
box 1986 -3967 2714 388
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_3 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform -1 0 147072 0 1 1458
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_5
timestamp 1715205430
transform -1 0 147072 0 1 6342
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_6
timestamp 1715205430
transform -1 0 147072 0 1 4714
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_7
timestamp 1715205430
transform -1 0 147072 0 1 3086
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_8
timestamp 1715205430
transform -1 0 144480 0 1 1458
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_9
timestamp 1715205430
transform -1 0 144480 0 1 4714
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_10
timestamp 1715205430
transform -1 0 144480 0 1 3086
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_11
timestamp 1715205430
transform -1 0 141888 0 1 1458
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_12
timestamp 1715205430
transform -1 0 144480 0 1 6342
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_13
timestamp 1715205430
transform -1 0 141888 0 1 6342
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_14
timestamp 1715205430
transform -1 0 141888 0 -1 3086
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_16
timestamp 1715205430
transform -1 0 141888 0 1 4714
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_17
timestamp 1715205430
transform -1 0 141888 0 1 3086
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_18
timestamp 1715205430
transform -1 0 141888 0 -1 4714
box -66 -43 450 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform -1 0 149280 0 -1 6342
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_1
timestamp 1715205430
transform -1 0 149280 0 -1 3086
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_2
timestamp 1715205430
transform -1 0 149280 0 -1 4714
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_3
timestamp 1715205430
transform -1 0 146688 0 1 1458
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_4
timestamp 1715205430
transform -1 0 149280 0 -1 7970
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_5
timestamp 1715205430
transform -1 0 146688 0 1 6342
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_6
timestamp 1715205430
transform -1 0 146688 0 1 4714
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_7
timestamp 1715205430
transform -1 0 146688 0 1 3086
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_8
timestamp 1715205430
transform -1 0 144096 0 1 1458
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_9
timestamp 1715205430
transform -1 0 144096 0 1 4714
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_10
timestamp 1715205430
transform -1 0 144096 0 1 3086
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_11
timestamp 1715205430
transform -1 0 141504 0 1 1458
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_12
timestamp 1715205430
transform -1 0 144096 0 1 6342
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_13
timestamp 1715205430
transform -1 0 141504 0 1 6342
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_14
timestamp 1715205430
transform -1 0 141504 0 -1 3086
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_16
timestamp 1715205430
transform -1 0 141504 0 1 4714
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_17
timestamp 1715205430
transform -1 0 141504 0 1 3086
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_18
timestamp 1715205430
transform -1 0 141504 0 -1 4714
box -66 -43 162 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform -1 0 147072 0 -1 3086
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_1
timestamp 1715205430
transform -1 0 141888 0 -1 7970
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_5
timestamp 1715205430
transform -1 0 147072 0 -1 7970
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_6
timestamp 1715205430
transform -1 0 147072 0 -1 6342
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_7
timestamp 1715205430
transform -1 0 147072 0 -1 4714
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_8
timestamp 1715205430
transform -1 0 144480 0 -1 4714
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_9
timestamp 1715205430
transform -1 0 144480 0 -1 3086
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_10
timestamp 1715205430
transform -1 0 144480 0 -1 7970
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_11
timestamp 1715205430
transform -1 0 144480 0 -1 6342
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_12
timestamp 1715205430
transform -1 0 141888 0 -1 6342
box -66 -43 546 897
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
array 0 3 -2592 0 3 1628
timestamp 1715205430
transform -1 0 141408 0 1 1458
box -66 -43 2178 1671
<< labels >>
flabel metal4 148877 1311 149477 2511 0 FreeSans 3200 90 0 0 dvss
port 4 nsew
flabel metal4 148877 2799 149477 4484 0 FreeSans 3200 90 0 0 avss
port 2 nsew
flabel metal4 66 2799 299 4484 0 FreeSans 1600 90 0 0 avss
port 2 nsew
flabel metal4 148877 4635 149477 6320 0 FreeSans 3200 90 0 0 avdd
port 1 nsew
flabel metal4 65 4635 298 6320 0 FreeSans 1600 90 0 0 avdd
port 1 nsew
flabel metal4 148877 6683 149477 7883 0 FreeSans 3200 90 0 0 dvdd
port 3 nsew
flabel metal3 136670 193 136875 335 0 FreeSans 1600 90 0 0 snk_test1
port 4 nsew
flabel metal3 136664 9225 136907 9466 0 FreeSans 1600 90 0 0 src_test1
port 5 nsew
flabel metal3 135980 9225 136219 9465 0 FreeSans 1600 90 0 0 src_50
port 6 nsew
flabel metal3 135551 9225 135909 9465 0 FreeSans 1600 90 0 0 src_100
port 7 nsew
flabel metal3 133999 9225 134357 9465 0 FreeSans 1600 90 0 0 src_200_2
port 8 nsew
flabel metal3 131907 9225 132265 9465 0 FreeSans 1600 90 0 0 src_200_1
port 9 nsew
flabel metal3 129815 9225 130173 9465 0 FreeSans 1600 90 0 0 src_200_0
port 10 nsew
flabel metal3 126645 9225 127003 9465 0 FreeSans 1600 90 0 0 src_400
port 11 nsew
flabel metal3 121385 9224 121747 9465 0 FreeSans 1600 90 0 0 src_600
port 12 nsew
flabel metal3 41543 9224 41905 9465 0 FreeSans 1600 90 0 0 src_10000
port 13 nsew
flabel metal3 137060 195 137194 337 0 FreeSans 1600 90 0 0 ena_test1_3v3
flabel metal3 137011 9226 137210 9467 0 FreeSans 1600 90 0 0 enb_test1_3v3
flabel metal3 136322 9225 136543 9465 0 FreeSans 1600 90 0 0 enb_50_3v3
flabel metal3 135196 9225 135417 9465 0 FreeSans 1600 90 0 0 enb_100_3v3
flabel metal3 133104 9225 133325 9465 0 FreeSans 1600 90 0 0 enb_200_2_3v3
flabel metal3 131012 9225 131233 9465 0 FreeSans 1600 90 0 0 enb_200_1_3v3
flabel metal3 128920 9225 129141 9465 0 FreeSans 1600 90 0 0 enb_200_0_3v3
flabel metal3 125750 9225 125971 9465 0 FreeSans 1600 90 0 0 enb_400_3v3
flabel metal3 120490 9225 120711 9466 0 FreeSans 1600 90 0 0 enb_600_3v3
flabel metal3 40664 9250 40885 9465 0 FreeSans 1600 90 0 0 enb_10000_3v3
flabel metal3 105479 1 105700 230 0 FreeSans 1600 90 0 0 ena_2000_3v3
flabel metal3 85706 0 85927 229 0 FreeSans 1600 90 0 0 ena_4000_3v3
flabel metal3 36199 0 36420 229 0 FreeSans 1600 90 0 0 ena_5000_3v3
flabel metal3 119987 1 120208 189 0 FreeSans 1600 90 0 0 ena_1000_3v3
flabel metal3 135060 195 135194 337 0 FreeSans 1600 90 0 0 ena_750_3v3
flabel metal3 111922 9224 112143 9465 0 FreeSans 1600 90 0 0 enb_1000_3v3
flabel metal3 120882 1 121244 189 0 FreeSans 1600 90 0 0 snk_1000
port 14 nsew
flabel metal3 134670 193 134875 335 0 FreeSans 1600 90 0 0 snk_750
port 15 nsew
flabel metal3 112817 9224 113179 9465 0 FreeSans 1600 90 0 0 src_1000
port 16 nsew
flabel metal3 106374 1 106736 230 0 FreeSans 1600 90 0 0 snk_2000
port 17 nsew
flabel metal3 86601 0 86963 229 0 FreeSans 1600 90 0 0 snk_4000
port 18 nsew
flabel metal3 37094 0 37456 229 0 FreeSans 1600 90 0 0 snk_5000
port 19 nsew
flabel metal2 143631 678 143671 1078 0 FreeSans 400 90 0 0 ena_snk_test1
port 20 nsew
flabel metal2 143751 678 143791 1053 0 FreeSans 400 90 0 0 ena_snk_750
port 21 nsew
flabel metal2 141039 678 141079 1053 0 FreeSans 400 90 0 0 ena_snk_1000
port 22 nsew
flabel metal2 141159 678 141199 1053 0 FreeSans 400 90 0 0 ena_snk_2000
port 23 nsew
flabel metal2 141279 678 141319 1053 0 FreeSans 400 90 0 0 ena_snk_4000
port 24 nsew
flabel metal2 141399 678 141439 1053 0 FreeSans 400 90 0 0 ena_snk_5000
port 25 nsew
flabel metal2 143991 678 144031 1053 0 FreeSans 400 90 0 0 ena_src_test1
port 26 nsew
flabel metal2 143871 678 143911 1053 0 FreeSans 400 90 0 0 ena_src_50
port 27 nsew
flabel metal2 146463 678 146503 1053 0 FreeSans 400 90 0 0 ena_src_100
port 28 nsew
flabel metal2 146583 678 146623 1053 0 FreeSans 400 90 0 0 ena_src_200_2
port 29 nsew
flabel metal2 146343 678 146383 1053 0 FreeSans 400 90 0 0 ena_src_200_1
port 30 nsew
flabel metal2 146223 678 146263 1053 0 FreeSans 400 90 0 0 ena_src_200_0
port 31 nsew
flabel metal2 149055 678 149095 1053 0 FreeSans 400 90 0 0 ena_src_400
port 32 nsew
flabel metal2 149175 678 149215 1053 0 FreeSans 400 90 0 0 ena_src_600
port 33 nsew
flabel metal2 148935 678 148975 1053 0 FreeSans 400 90 0 0 ena_src_1000
port 34 nsew
flabel metal2 148815 678 148855 1053 0 FreeSans 400 90 0 0 ena_src_10000
port 35 nsew
<< end >>
