magic
tech sky130A
magscale 1 2
timestamp 1716927123
<< error_s >>
rect 66 8804 90 8828
rect 42 8770 66 8804
rect 66 8746 90 8770
rect 0 8618 66 8680
rect 0 8614 90 8618
rect 0 8540 132 8614
rect 0 8536 90 8540
rect 0 8474 66 8536
rect 66 925 966 1825
rect 0 754 66 816
rect 0 750 90 754
rect 0 676 132 750
rect 0 672 90 676
rect 0 610 66 672
rect 66 522 72 523
rect 66 498 90 522
rect 42 479 72 498
rect 42 464 66 479
rect 66 440 90 464
<< dnwell >>
rect 66 719 138229 8571
<< nwell >>
rect 66 8365 138338 8680
rect 138023 925 138338 8365
rect 66 610 138338 925
<< pwell >>
rect 2095 925 2183 947
<< mvpsubdiff >>
rect 138398 8770 138458 8804
rect 138424 8744 138458 8770
rect 139072 8182 139132 8216
rect 149416 8182 149476 8216
rect 139072 8156 139106 8182
rect 139072 1252 139106 1278
rect 149442 8156 149476 8182
rect 149442 1252 149476 1278
rect 139072 1218 139132 1252
rect 149416 1218 149476 1252
rect 138424 498 138458 524
rect 138398 464 138458 498
<< mvnsubdiff >>
rect 66 8594 138272 8614
rect 138192 8560 138272 8594
rect 66 8540 138272 8560
rect 138198 8534 138272 8540
rect 138198 756 138218 8534
rect 138252 756 138272 8534
rect 138198 750 138272 756
rect 66 730 138272 750
rect 138192 696 138272 730
rect 66 676 138272 696
<< mvpsubdiffcont >>
rect 66 8770 138398 8804
rect 138424 524 138458 8744
rect 139132 8182 149416 8216
rect 139072 1278 139106 8156
rect 149442 1278 149476 8156
rect 139132 1218 149416 1252
rect 66 464 138398 498
<< mvnsubdiffcont >>
rect 66 8560 138192 8594
rect 138218 756 138252 8534
rect 66 696 138192 730
<< locali >>
rect 138398 8770 138458 8804
rect 66 8755 138458 8770
rect 66 8671 138360 8755
rect 138192 8560 138252 8594
rect 66 8534 138252 8560
rect 66 8529 138218 8534
rect 66 8375 138128 8529
rect 138081 909 138128 8375
rect 66 752 138128 909
rect 138187 756 138218 8529
rect 138187 752 138252 756
rect 66 730 138252 752
rect 138192 696 138252 730
rect 138316 610 138360 8671
rect 66 523 138360 610
rect 138307 514 138360 523
rect 138412 8744 138458 8755
rect 138412 524 138424 8744
rect 139072 8182 139132 8216
rect 149416 8182 149476 8216
rect 139072 8156 149476 8182
rect 139106 8094 149442 8156
rect 139106 1340 139189 8094
rect 141863 7594 141910 7660
rect 144455 7594 144502 7660
rect 147047 7594 147094 7660
rect 140909 6766 141079 6782
rect 140909 6664 140925 6766
rect 141058 6664 141079 6766
rect 140909 6648 141079 6664
rect 143501 6766 143671 6782
rect 143501 6664 143517 6766
rect 143650 6664 143671 6766
rect 143501 6648 143671 6664
rect 146093 6766 146263 6782
rect 146093 6664 146109 6766
rect 146242 6664 146263 6766
rect 146093 6648 146263 6664
rect 148685 6766 148855 6782
rect 148685 6664 148701 6766
rect 148834 6664 148855 6766
rect 148685 6648 148855 6664
rect 141863 5966 141910 6032
rect 144455 5966 144502 6032
rect 147047 5966 147094 6032
rect 140909 5138 141079 5154
rect 140909 5036 140925 5138
rect 141058 5036 141079 5138
rect 140909 5020 141079 5036
rect 143501 5138 143671 5154
rect 143501 5036 143517 5138
rect 143650 5036 143671 5138
rect 143501 5020 143671 5036
rect 146093 5138 146263 5154
rect 146093 5036 146109 5138
rect 146242 5036 146263 5138
rect 146093 5020 146263 5036
rect 148685 5138 148855 5154
rect 148685 5036 148701 5138
rect 148834 5036 148855 5138
rect 148685 5020 148855 5036
rect 144455 4338 144502 4404
rect 147047 4338 147094 4404
rect 140909 3510 141079 3526
rect 140909 3408 140925 3510
rect 141058 3408 141079 3510
rect 140909 3392 141079 3408
rect 143501 3510 143671 3526
rect 143501 3408 143517 3510
rect 143650 3408 143671 3510
rect 143501 3392 143671 3408
rect 146093 3510 146263 3526
rect 146093 3408 146109 3510
rect 146242 3408 146263 3510
rect 146093 3392 146263 3408
rect 148685 3510 148855 3526
rect 148685 3408 148701 3510
rect 148834 3408 148855 3510
rect 148685 3392 148855 3408
rect 144455 2710 144502 2776
rect 147047 2710 147094 2776
rect 140909 1882 141079 1898
rect 140909 1780 140925 1882
rect 141058 1780 141079 1882
rect 140909 1764 141079 1780
rect 143501 1882 143671 1898
rect 143501 1780 143517 1882
rect 143650 1780 143671 1882
rect 143501 1764 143671 1780
rect 146093 1882 146263 1898
rect 146093 1780 146109 1882
rect 146242 1780 146263 1882
rect 146093 1764 146263 1780
rect 148685 1882 148855 1898
rect 148685 1780 148701 1882
rect 148834 1780 148855 1882
rect 148685 1764 148855 1780
rect 149348 1340 149442 8094
rect 139106 1278 149442 1340
rect 139072 1252 149476 1278
rect 139072 1218 139132 1252
rect 149416 1218 149476 1252
rect 138412 514 138458 524
rect 138307 498 138458 514
rect 138398 464 138458 498
<< viali >>
rect 138128 752 138187 8529
rect 66 498 138307 523
rect 138360 514 138412 8755
rect 141529 7624 141575 7803
rect 144121 7624 144167 7803
rect 146713 7624 146759 7803
rect 139318 7316 139366 7547
rect 140925 6664 141058 6766
rect 143517 6664 143650 6766
rect 146109 6664 146242 6766
rect 148701 6664 148834 6766
rect 141529 5996 141575 6175
rect 144121 5996 144167 6175
rect 146713 5996 146759 6175
rect 139318 5688 139366 5919
rect 140925 5036 141058 5138
rect 143517 5036 143650 5138
rect 146109 5036 146242 5138
rect 148701 5036 148834 5138
rect 144121 4368 144167 4547
rect 146713 4368 146759 4547
rect 139318 4060 139366 4291
rect 141910 4060 141958 4291
rect 140925 3408 141058 3510
rect 143517 3408 143650 3510
rect 146109 3408 146242 3510
rect 148701 3408 148834 3510
rect 144121 2740 144167 2919
rect 146713 2740 146759 2919
rect 139318 2432 139366 2663
rect 141910 2432 141958 2663
rect 140925 1780 141058 1882
rect 143517 1780 143650 1882
rect 146109 1780 146242 1882
rect 148701 1780 148834 1882
rect 66 479 138307 498
<< metal1 >>
rect 138332 8755 138448 8797
rect 138093 8529 138231 8580
rect 138093 6299 138128 8529
rect 138187 6299 138231 8529
rect 33780 5926 33848 6035
rect 33630 5692 33780 5894
rect 33630 5648 33848 5692
rect 138093 4657 138108 6299
rect 138215 4657 138231 6299
rect 23115 3456 23177 3471
rect 23115 3125 23177 3218
rect 23649 3456 23711 3471
rect 23649 3125 23711 3218
rect 24183 3456 24245 3471
rect 24183 3125 24245 3218
rect 24717 3456 24779 3471
rect 24717 3125 24779 3218
rect 25251 3456 25313 3471
rect 25251 3125 25313 3218
rect 25785 3456 25847 3471
rect 25785 3125 25847 3218
rect 26319 3456 26381 3471
rect 26319 3125 26381 3218
rect 26853 3456 26915 3471
rect 26853 3125 26915 3218
rect 27387 3456 27449 3471
rect 27387 3125 27449 3218
rect 27921 3456 27983 3471
rect 27921 3125 27983 3218
rect 28455 3456 28517 3471
rect 28455 3125 28517 3218
rect 28989 3456 29051 3471
rect 28989 3125 29051 3218
rect 29523 3456 29585 3471
rect 29523 3125 29585 3218
rect 30057 3456 30119 3471
rect 30057 3125 30119 3218
rect 30591 3456 30653 3471
rect 30591 3125 30653 3218
rect 31125 3456 31187 3471
rect 31125 3125 31187 3218
rect 31659 3456 31721 3471
rect 31659 3125 31721 3218
rect 32193 3456 32255 3471
rect 32193 3125 32255 3218
rect 32727 3456 32789 3471
rect 32727 3125 32789 3218
rect 33261 3456 33323 3471
rect 33261 3125 33323 3218
rect 23315 2472 23379 2482
rect 23315 2159 23379 2234
rect 23849 2472 23913 2482
rect 23849 2159 23913 2234
rect 24383 2472 24447 2482
rect 24383 2159 24447 2234
rect 24917 2472 24981 2482
rect 24917 2159 24981 2234
rect 25451 2472 25515 2482
rect 25451 2159 25515 2234
rect 25985 2472 26049 2482
rect 25985 2159 26049 2234
rect 26511 2472 26583 2482
rect 26511 2159 26583 2234
rect 27045 2472 27117 2482
rect 27045 2159 27117 2234
rect 27579 2472 27651 2482
rect 27579 2159 27651 2234
rect 28113 2472 28185 2482
rect 28113 2159 28185 2234
rect 28647 2472 28719 2482
rect 28647 2159 28719 2234
rect 29181 2472 29253 2482
rect 29181 2159 29253 2234
rect 29715 2472 29787 2482
rect 29715 2159 29787 2234
rect 30249 2472 30321 2482
rect 30249 2159 30321 2234
rect 30783 2472 30847 2482
rect 30783 2159 30847 2234
rect 31317 2472 31381 2482
rect 31317 2159 31381 2234
rect 31851 2472 31915 2482
rect 31851 2159 31915 2234
rect 32385 2472 32449 2482
rect 32385 2159 32449 2234
rect 32919 2472 32983 2482
rect 32919 2159 32983 2234
rect 23489 821 23543 849
rect 24023 821 24077 849
rect 24557 821 24611 849
rect 25091 821 25145 849
rect 25625 821 25679 849
rect 26159 821 26213 849
rect 26693 821 26747 849
rect 27227 821 27281 849
rect 27761 821 27815 849
rect 28295 821 28349 849
rect 28829 821 28883 849
rect 29363 821 29417 849
rect 29897 821 29951 849
rect 30431 821 30485 849
rect 30965 821 31019 849
rect 31499 821 31553 849
rect 32033 821 32087 849
rect 32567 821 32621 849
rect 33101 821 33155 849
rect 33635 821 33689 849
rect 138093 752 138128 4657
rect 138187 752 138231 4657
rect 138093 705 138231 752
rect 138332 542 138360 8755
rect 66 523 138360 542
rect 138307 514 138360 523
rect 138412 514 138448 8755
rect 141522 7803 141581 7815
rect 141522 7784 141529 7803
rect 139006 7744 141529 7784
rect 139006 7664 141400 7704
rect 139006 7584 141296 7624
rect 139306 7547 139384 7553
rect 139306 7544 139318 7547
rect 139006 7504 139318 7544
rect 139306 7316 139318 7504
rect 139366 7316 139384 7547
rect 141256 7442 141296 7584
rect 141360 7529 141400 7664
rect 141522 7624 141529 7744
rect 141575 7624 141581 7803
rect 141522 7612 141581 7624
rect 144114 7803 144173 7815
rect 144114 7624 144121 7803
rect 144167 7624 144173 7803
rect 144114 7612 144173 7624
rect 146706 7803 146765 7815
rect 146706 7624 146713 7803
rect 146759 7624 146765 7803
rect 146706 7612 146765 7624
rect 144132 7529 144172 7612
rect 141360 7489 144172 7529
rect 146720 7442 146760 7612
rect 141256 7402 146760 7442
rect 139306 7310 139384 7316
rect 140909 6766 141079 6782
rect 140909 6664 140925 6766
rect 141058 6664 141079 6766
rect 140909 6648 141079 6664
rect 143501 6766 143671 6782
rect 143501 6664 143517 6766
rect 143650 6664 143671 6766
rect 143501 6648 143671 6664
rect 146093 6766 146263 6782
rect 146093 6664 146109 6766
rect 146242 6664 146263 6766
rect 146093 6648 146263 6664
rect 148685 6766 148855 6782
rect 148685 6664 148701 6766
rect 148834 6664 148855 6766
rect 148685 6648 148855 6664
rect 141522 6175 141581 6187
rect 141522 6156 141529 6175
rect 139006 6116 141529 6156
rect 139006 6036 141400 6076
rect 139006 5956 141296 5996
rect 139306 5919 139384 5925
rect 139306 5916 139318 5919
rect 139006 5876 139318 5916
rect 139306 5688 139318 5876
rect 139366 5688 139384 5919
rect 141256 5814 141296 5956
rect 141360 5901 141400 6036
rect 141522 5996 141529 6116
rect 141575 5996 141581 6175
rect 141522 5984 141581 5996
rect 144114 6175 144173 6187
rect 144114 5996 144121 6175
rect 144167 5996 144173 6175
rect 144114 5984 144173 5996
rect 146706 6175 146765 6187
rect 146706 5996 146713 6175
rect 146759 5996 146765 6175
rect 146706 5984 146765 5996
rect 144132 5901 144172 5984
rect 141360 5861 144172 5901
rect 146720 5814 146760 5984
rect 141256 5774 146760 5814
rect 139306 5682 139384 5688
rect 140909 5138 141079 5154
rect 140909 5036 140925 5138
rect 141058 5036 141079 5138
rect 140909 5020 141079 5036
rect 143501 5138 143671 5154
rect 143501 5036 143517 5138
rect 143650 5036 143671 5138
rect 143501 5020 143671 5036
rect 146093 5138 146263 5154
rect 146093 5036 146109 5138
rect 146242 5036 146263 5138
rect 146093 5020 146263 5036
rect 148685 5138 148855 5154
rect 148685 5036 148701 5138
rect 148834 5036 148855 5138
rect 148685 5020 148855 5036
rect 144114 4547 144173 4559
rect 144114 4528 144121 4547
rect 139006 4488 144121 4528
rect 139006 4408 143157 4448
rect 139006 4328 141959 4368
rect 141919 4297 141959 4328
rect 139306 4291 139384 4297
rect 139306 4288 139318 4291
rect 139006 4248 139318 4288
rect 139306 4060 139318 4248
rect 139366 4060 139384 4291
rect 139306 4054 139384 4060
rect 141898 4291 141976 4297
rect 141898 4060 141910 4291
rect 141958 4060 141976 4291
rect 143117 4186 143157 4408
rect 144114 4368 144121 4488
rect 144167 4368 144173 4547
rect 144114 4356 144173 4368
rect 146706 4547 146765 4559
rect 146706 4368 146713 4547
rect 146759 4368 146765 4547
rect 146706 4356 146765 4368
rect 146720 4186 146760 4356
rect 143117 4146 146760 4186
rect 141898 4054 141976 4060
rect 140909 3510 141079 3526
rect 140909 3408 140925 3510
rect 141058 3408 141079 3510
rect 140909 3392 141079 3408
rect 143501 3510 143671 3526
rect 143501 3408 143517 3510
rect 143650 3408 143671 3510
rect 143501 3392 143671 3408
rect 146093 3510 146263 3526
rect 146093 3408 146109 3510
rect 146242 3408 146263 3510
rect 146093 3392 146263 3408
rect 148685 3510 148855 3526
rect 148685 3408 148701 3510
rect 148834 3408 148855 3510
rect 148685 3392 148855 3408
rect 144114 2919 144173 2931
rect 144114 2900 144121 2919
rect 139006 2860 144121 2900
rect 139006 2780 143208 2820
rect 139006 2700 141955 2740
rect 141915 2669 141955 2700
rect 139306 2663 139384 2669
rect 139306 2660 139318 2663
rect 139006 2620 139318 2660
rect 139306 2432 139318 2620
rect 139366 2432 139384 2663
rect 139306 2426 139384 2432
rect 141898 2663 141976 2669
rect 141898 2432 141910 2663
rect 141958 2432 141976 2663
rect 143168 2558 143208 2780
rect 144114 2740 144121 2860
rect 144167 2740 144173 2919
rect 144114 2728 144173 2740
rect 146706 2919 146765 2931
rect 146706 2740 146713 2919
rect 146759 2740 146765 2919
rect 146706 2728 146765 2740
rect 146720 2558 146760 2728
rect 143168 2518 146760 2558
rect 141898 2426 141976 2432
rect 140909 1882 141079 1898
rect 140909 1780 140925 1882
rect 141058 1780 141079 1882
rect 140909 1764 141079 1780
rect 143501 1882 143671 1898
rect 143501 1780 143517 1882
rect 143650 1780 143671 1882
rect 143501 1764 143671 1780
rect 146093 1882 146263 1898
rect 146093 1780 146109 1882
rect 146242 1780 146263 1882
rect 146093 1764 146263 1780
rect 148685 1882 148855 1898
rect 148685 1780 148701 1882
rect 148834 1780 148855 1882
rect 148685 1764 148855 1780
rect 138307 479 138448 514
rect 66 464 138448 479
<< via1 >>
rect 33634 8737 33688 8969
rect 33475 7030 33544 7589
rect 33780 5692 33848 5926
rect 138108 4657 138128 6299
rect 138128 4657 138187 6299
rect 138187 4657 138215 6299
rect 23115 3218 23177 3456
rect 23649 3218 23711 3456
rect 24183 3218 24245 3456
rect 24717 3218 24779 3456
rect 25251 3218 25313 3456
rect 25785 3218 25847 3456
rect 26319 3218 26381 3456
rect 26853 3218 26915 3456
rect 27387 3218 27449 3456
rect 27921 3218 27983 3456
rect 28455 3218 28517 3456
rect 28989 3218 29051 3456
rect 29523 3218 29585 3456
rect 30057 3218 30119 3456
rect 30591 3218 30653 3456
rect 31125 3218 31187 3456
rect 31659 3218 31721 3456
rect 32193 3218 32255 3456
rect 32727 3218 32789 3456
rect 33261 3218 33323 3456
rect 23315 2234 23379 2472
rect 23849 2234 23913 2472
rect 24383 2234 24447 2472
rect 24917 2234 24981 2472
rect 25451 2234 25515 2472
rect 25985 2234 26049 2472
rect 26511 2234 26583 2472
rect 27045 2234 27117 2472
rect 27579 2234 27651 2472
rect 28113 2234 28185 2472
rect 28647 2234 28719 2472
rect 29181 2234 29253 2472
rect 29715 2234 29787 2472
rect 30249 2234 30321 2472
rect 30783 2234 30847 2472
rect 31317 2234 31381 2472
rect 31851 2234 31915 2472
rect 32385 2234 32449 2472
rect 32919 2234 32983 2472
rect 33469 1579 33557 2146
rect 23489 849 23543 1037
rect 24023 849 24077 1037
rect 24557 849 24611 1037
rect 25091 849 25145 1037
rect 25625 849 25679 1037
rect 26159 849 26213 1037
rect 26693 849 26747 1037
rect 27227 849 27281 1037
rect 27761 849 27815 1037
rect 28295 849 28349 1037
rect 28829 849 28883 1037
rect 29363 849 29417 1037
rect 29897 849 29951 1037
rect 30431 849 30485 1037
rect 30965 849 31019 1037
rect 31499 849 31553 1037
rect 32033 849 32087 1037
rect 32567 849 32621 1037
rect 33101 849 33155 1037
rect 33635 849 33689 1037
rect 140925 6664 141058 6766
rect 143517 6664 143650 6766
rect 146109 6664 146242 6766
rect 148701 6664 148834 6766
rect 140925 5036 141058 5138
rect 143517 5036 143650 5138
rect 146109 5036 146242 5138
rect 148701 5036 148834 5138
rect 140925 3408 141058 3510
rect 143517 3408 143650 3510
rect 146109 3408 146242 3510
rect 148701 3408 148834 3510
rect 140925 1780 141058 1882
rect 143517 1780 143650 1882
rect 146109 1780 146242 1882
rect 148701 1780 148834 1882
<< metal2 >>
rect 33557 8969 33725 9237
rect 331 8735 33290 8967
rect 33376 8735 33385 8967
rect 33557 8737 33634 8969
rect 33688 8737 33725 8969
rect 517 8428 33292 8660
rect 33378 8428 33389 8660
rect 33557 8418 33725 8737
rect 33762 8735 33772 8967
rect 33858 8735 41568 8967
rect 41887 8735 54234 8967
rect 54561 8735 117480 8967
rect 117754 8735 121402 8967
rect 121729 8735 123820 8967
rect 124170 8735 126662 8967
rect 126989 8735 128250 8967
rect 128539 8735 129832 8967
rect 130159 8735 130497 8967
rect 130685 8735 131924 8967
rect 132251 8735 132590 8967
rect 132825 8735 134016 8967
rect 134343 8735 134797 8967
rect 134929 8735 135568 8967
rect 135895 8735 135909 8967
rect 135981 8735 135997 8967
rect 136169 8735 136203 8967
rect 136506 8735 136678 8967
rect 136895 8735 137113 8967
rect 33761 8428 33772 8660
rect 33858 8428 40683 8660
rect 40866 8428 53339 8660
rect 53524 8428 117627 8660
rect 117926 8428 120507 8660
rect 120692 8428 123968 8660
rect 124197 8428 125767 8660
rect 125952 8428 128328 8660
rect 128617 8428 128937 8660
rect 129122 8428 130589 8660
rect 130721 8428 131029 8660
rect 131214 8428 132590 8660
rect 132825 8428 133121 8660
rect 133306 8428 134797 8660
rect 134929 8428 135213 8660
rect 135398 8428 135858 8660
rect 135981 8428 136339 8660
rect 136524 8428 136549 8660
rect 136693 8428 137022 8660
rect 137197 8428 137292 8660
rect 66 8027 137616 8265
rect 66 7696 188 7930
rect 137608 7696 137655 7930
rect 137910 7696 137939 7930
rect 33475 7589 33544 7598
rect 33475 7021 33544 7030
rect 66 6696 137616 6930
rect 140909 6766 141079 6782
rect 66 6695 186 6696
rect 140909 6664 140925 6766
rect 141058 6739 141079 6766
rect 143501 6766 143671 6782
rect 141058 6699 141439 6739
rect 141058 6664 141079 6699
rect 140909 6648 141079 6664
rect 138079 6299 138248 6321
rect 182 5692 33780 5926
rect 33848 5692 137616 5926
rect 137608 4638 137654 4872
rect 137909 4638 137938 4872
rect 138079 4657 138108 6299
rect 138215 4657 138248 6299
rect 140909 5138 141079 5154
rect 140909 5036 140925 5138
rect 141058 5097 141079 5138
rect 141058 5057 141319 5097
rect 141058 5036 141079 5057
rect 140909 5020 141079 5036
rect 138079 4638 138248 4657
rect 66 4461 1279 4480
rect 66 4377 318 4461
rect 66 4242 1279 4377
rect 140909 3510 141079 3526
rect 223 3218 23115 3456
rect 23177 3218 23649 3456
rect 23711 3218 24183 3456
rect 24245 3218 24717 3456
rect 24779 3218 25251 3456
rect 25313 3218 25785 3456
rect 25847 3218 26319 3456
rect 26381 3218 26853 3456
rect 26915 3218 27387 3456
rect 27449 3218 27921 3456
rect 27983 3218 28455 3456
rect 28517 3218 28989 3456
rect 29051 3218 29523 3456
rect 29585 3218 30057 3456
rect 30119 3218 30591 3456
rect 30653 3218 31125 3456
rect 31187 3218 31659 3456
rect 31721 3218 32193 3456
rect 32255 3218 32727 3456
rect 32789 3218 33261 3456
rect 33323 3218 137597 3456
rect 140909 3408 140925 3510
rect 141058 3474 141079 3510
rect 141058 3434 141199 3474
rect 141058 3408 141079 3434
rect 140909 3392 141079 3408
rect 165 2234 23315 2472
rect 23379 2234 23849 2472
rect 23913 2234 24383 2472
rect 24447 2234 24917 2472
rect 24981 2234 25451 2472
rect 25515 2234 25985 2472
rect 26049 2234 26511 2472
rect 26583 2234 27045 2472
rect 27117 2234 27579 2472
rect 27651 2234 28113 2472
rect 28185 2234 28647 2472
rect 28719 2234 29181 2472
rect 29253 2234 29715 2472
rect 29787 2234 30249 2472
rect 30321 2234 30783 2472
rect 30847 2234 31317 2472
rect 31381 2234 31851 2472
rect 31915 2234 32385 2472
rect 32449 2234 32919 2472
rect 32983 2234 137589 2472
rect 33469 2146 33557 2155
rect 140909 1882 141079 1898
rect 140909 1780 140925 1882
rect 141058 1780 141079 1882
rect 140909 1764 141079 1780
rect 33469 1570 33557 1579
rect 66 1246 137597 1484
rect 141039 1134 141079 1764
rect 141159 1134 141199 3434
rect 141279 1134 141319 5057
rect 141399 1134 141439 6699
rect 143501 6664 143517 6766
rect 143650 6739 143671 6766
rect 146093 6766 146263 6782
rect 143650 6699 144031 6739
rect 143650 6664 143671 6699
rect 143501 6648 143671 6664
rect 143501 5138 143671 5154
rect 143501 5036 143517 5138
rect 143650 5097 143671 5138
rect 143650 5057 143911 5097
rect 143650 5036 143671 5057
rect 143501 5020 143671 5036
rect 143501 3510 143671 3526
rect 143501 3408 143517 3510
rect 143650 3474 143671 3510
rect 143650 3434 143791 3474
rect 143650 3408 143671 3434
rect 143501 3392 143671 3408
rect 143501 1882 143671 1898
rect 143501 1780 143517 1882
rect 143650 1780 143671 1882
rect 143501 1764 143671 1780
rect 143631 1134 143671 1764
rect 143751 1134 143791 3434
rect 143871 1134 143911 5057
rect 143991 1134 144031 6699
rect 146093 6664 146109 6766
rect 146242 6739 146263 6766
rect 148685 6766 148855 6782
rect 146242 6699 146623 6739
rect 146242 6664 146263 6699
rect 146093 6648 146263 6664
rect 146093 5138 146263 5154
rect 146093 5036 146109 5138
rect 146242 5097 146263 5138
rect 146242 5057 146503 5097
rect 146242 5036 146263 5057
rect 146093 5020 146263 5036
rect 146093 3510 146263 3526
rect 146093 3408 146109 3510
rect 146242 3474 146263 3510
rect 146242 3434 146383 3474
rect 146242 3408 146263 3434
rect 146093 3392 146263 3408
rect 146093 1882 146263 1898
rect 146093 1780 146109 1882
rect 146242 1780 146263 1882
rect 146093 1764 146263 1780
rect 146223 1134 146263 1764
rect 146343 1134 146383 3434
rect 146463 1134 146503 5057
rect 146583 1134 146623 6699
rect 148685 6664 148701 6766
rect 148834 6739 148855 6766
rect 148834 6699 149215 6739
rect 148834 6664 148855 6699
rect 148685 6648 148855 6664
rect 148685 5138 148855 5154
rect 148685 5036 148701 5138
rect 148834 5097 148855 5138
rect 148834 5057 149095 5097
rect 148834 5036 148855 5057
rect 148685 5020 148855 5036
rect 148685 3510 148855 3526
rect 148685 3408 148701 3510
rect 148834 3474 148855 3510
rect 148834 3434 148975 3474
rect 148834 3408 148855 3434
rect 148685 3392 148855 3408
rect 148685 1882 148855 1898
rect 148685 1780 148701 1882
rect 148834 1780 148855 1882
rect 148685 1764 148855 1780
rect 148815 1134 148855 1764
rect 148935 1134 148975 3434
rect 149055 1134 149095 5057
rect 149175 1134 149215 6699
rect 66 849 10216 1037
rect 10401 849 22503 1037
rect 22567 849 23489 1037
rect 23543 849 24023 1037
rect 24077 849 24557 1037
rect 24611 849 25091 1037
rect 25145 849 25625 1037
rect 25679 849 26159 1037
rect 26213 849 26693 1037
rect 26747 849 27227 1037
rect 27281 849 27761 1037
rect 27815 849 28295 1037
rect 28349 849 28829 1037
rect 28883 849 29363 1037
rect 29417 849 29897 1037
rect 29951 849 30431 1037
rect 30485 849 30965 1037
rect 31019 849 31499 1037
rect 31553 849 32033 1037
rect 32087 849 32567 1037
rect 32621 849 33101 1037
rect 33155 849 33635 1037
rect 33689 849 33855 1037
rect 34152 849 63896 1037
rect 64081 849 96188 1037
rect 96610 849 120004 1037
rect 120189 849 136239 1037
rect 136690 849 137068 1037
rect 137185 849 137300 1037
rect 66 593 11111 781
rect 11438 593 22335 781
rect 22567 763 22667 849
rect 22467 563 22667 763
rect 22753 593 32999 781
rect 33431 593 33523 781
rect 33981 593 64791 781
rect 65118 593 96022 781
rect 96444 593 120899 781
rect 121226 593 136081 781
rect 136525 593 136680 781
rect 136862 593 137135 781
<< via2 >>
rect 33290 8735 33376 8967
rect 33292 8428 33378 8660
rect 33772 8735 33858 8967
rect 41568 8735 41887 8967
rect 54234 8735 54561 8967
rect 121402 8735 121729 8967
rect 126662 8735 126989 8967
rect 129832 8735 130159 8967
rect 131924 8735 132251 8967
rect 134016 8735 134343 8967
rect 135568 8735 135895 8967
rect 135997 8735 136169 8967
rect 136678 8735 136895 8967
rect 33772 8428 33858 8660
rect 40683 8428 40866 8660
rect 53339 8428 53524 8660
rect 120507 8428 120692 8660
rect 125767 8428 125952 8660
rect 128937 8428 129122 8660
rect 131029 8428 131214 8660
rect 133121 8428 133306 8660
rect 135213 8428 135398 8660
rect 136339 8428 136524 8660
rect 137022 8428 137197 8660
rect 137655 7696 137910 7930
rect 33475 7030 33544 7589
rect 317 4654 33298 4738
rect 33715 4654 137146 4738
rect 137654 4638 137909 4872
rect 138108 4657 138215 6299
rect 318 4377 33299 4461
rect 33716 4379 137147 4463
rect 33469 1579 33557 2146
rect 10216 849 10401 1037
rect 63896 849 64081 1037
rect 120004 849 120189 1037
rect 137068 849 137185 1037
rect 11111 593 11438 781
rect 64791 593 65118 781
rect 120899 593 121226 781
rect 136680 593 136862 781
<< metal3 >>
rect 33284 8967 33866 8975
rect 33284 8735 33290 8967
rect 33376 8735 33772 8967
rect 33858 8735 33866 8967
rect 33284 8730 33866 8735
rect 33283 8660 33867 8668
rect 33283 8428 33292 8660
rect 33378 8428 33772 8660
rect 33858 8428 33867 8660
rect 33283 8418 33867 8428
rect 40664 8660 40885 9465
rect 41542 8967 41905 9465
rect 41542 8735 41568 8967
rect 41887 8735 41905 8967
rect 41542 8714 41905 8735
rect 40664 8428 40683 8660
rect 40866 8428 40885 8660
rect 40664 8390 40885 8428
rect 53322 8660 53543 9465
rect 54217 8967 54579 9465
rect 54217 8735 54234 8967
rect 54561 8735 54579 8967
rect 54217 8714 54579 8735
rect 53322 8428 53339 8660
rect 53524 8428 53543 8660
rect 53322 8390 53543 8428
rect 120490 8660 120711 9466
rect 121385 8967 121747 9465
rect 121385 8735 121402 8967
rect 121729 8735 121747 8967
rect 121385 8714 121747 8735
rect 120490 8428 120507 8660
rect 120692 8428 120711 8660
rect 120490 8390 120711 8428
rect 125750 8660 125971 9465
rect 126645 8967 127003 9465
rect 126645 8735 126662 8967
rect 126989 8735 127003 8967
rect 126645 8714 127003 8735
rect 125750 8428 125767 8660
rect 125952 8428 125971 8660
rect 125750 8390 125971 8428
rect 128920 8660 129141 9465
rect 129815 8967 130173 9465
rect 129815 8735 129832 8967
rect 130159 8735 130173 8967
rect 129815 8714 130173 8735
rect 128920 8428 128937 8660
rect 129122 8428 129141 8660
rect 128920 8390 129141 8428
rect 131012 8660 131233 9465
rect 131907 8967 132265 9465
rect 131907 8735 131924 8967
rect 132251 8735 132265 8967
rect 131907 8714 132265 8735
rect 131012 8428 131029 8660
rect 131214 8428 131233 8660
rect 131012 8390 131233 8428
rect 133104 8660 133325 9465
rect 133999 8967 134357 9465
rect 133999 8735 134016 8967
rect 134343 8735 134357 8967
rect 133999 8714 134357 8735
rect 133104 8428 133121 8660
rect 133306 8428 133325 8660
rect 133104 8390 133325 8428
rect 135196 8660 135417 9465
rect 135551 8967 135909 9465
rect 135551 8735 135568 8967
rect 135895 8735 135909 8967
rect 135551 8714 135909 8735
rect 135980 8967 136219 9465
rect 135980 8735 135997 8967
rect 136169 8735 136219 8967
rect 135980 8714 136219 8735
rect 135196 8428 135213 8660
rect 135398 8428 135417 8660
rect 135196 8390 135417 8428
rect 136322 8660 136543 9465
rect 136664 8967 136907 9466
rect 136664 8735 136678 8967
rect 136895 8735 136907 8967
rect 136664 8715 136907 8735
rect 136322 8428 136339 8660
rect 136524 8428 136543 8660
rect 136322 8390 136543 8428
rect 137011 8660 137210 9467
rect 137011 8428 137022 8660
rect 137197 8428 137210 8660
rect 137011 8408 137210 8428
rect 137642 7930 137920 7967
rect 137642 7696 137655 7930
rect 137910 7696 137920 7930
rect 33463 7589 33562 7657
rect 33463 7030 33475 7589
rect 33544 7030 33562 7589
rect 292 4827 33371 4872
rect 292 4654 317 4827
rect 33298 4654 33371 4827
rect 292 4638 33371 4654
rect 279 4461 33371 4480
rect 33299 4288 33371 4461
rect 279 4242 33371 4288
rect 33463 2146 33562 7030
rect 137642 4872 137920 7696
rect 33650 4827 137654 4872
rect 33650 4653 33715 4827
rect 137147 4653 137654 4827
rect 33650 4638 137654 4653
rect 137909 4638 137920 4872
rect 138079 6299 138248 6321
rect 138079 4657 138108 6299
rect 138215 4657 138248 6299
rect 138079 4638 138248 4657
rect 33650 4464 137539 4480
rect 33650 4290 33715 4464
rect 137147 4290 137539 4464
rect 33650 4242 137539 4290
rect 33463 1579 33469 2146
rect 33557 1579 33562 2146
rect 33463 1573 33562 1579
rect 137642 1254 137920 4638
rect 10199 1037 10420 1075
rect 10199 849 10216 1037
rect 10401 849 10420 1037
rect 10199 0 10420 849
rect 11094 781 11456 802
rect 11094 593 11111 781
rect 11438 593 11456 781
rect 11094 0 11456 593
rect 56506 0 56727 1075
rect 63879 1037 64100 1076
rect 63879 849 63896 1037
rect 64081 849 64100 1037
rect 57401 0 57763 802
rect 63879 1 64100 849
rect 119987 1037 120208 1076
rect 119987 849 120004 1037
rect 120189 849 120208 1037
rect 64774 781 65136 803
rect 64774 593 64791 781
rect 65118 593 65136 781
rect 64774 1 65136 593
rect 119987 1 120208 849
rect 137060 1037 137194 1053
rect 137060 849 137068 1037
rect 137185 849 137194 1037
rect 120882 781 121244 803
rect 120882 593 120899 781
rect 121226 593 121244 781
rect 120882 1 121244 593
rect 136670 781 136875 800
rect 136670 593 136680 781
rect 136862 593 136875 781
rect 136670 193 136875 593
rect 137060 195 137194 849
<< via3 >>
rect 317 4738 33298 4827
rect 317 4654 33298 4738
rect 279 4377 318 4461
rect 318 4377 33299 4461
rect 279 4288 33299 4377
rect 33715 4738 137147 4827
rect 33715 4654 137146 4738
rect 137146 4654 137147 4738
rect 33715 4653 137147 4654
rect 138108 4657 138215 6299
rect 33715 4463 137147 4464
rect 33715 4379 33716 4463
rect 33716 4379 137147 4463
rect 33715 4290 137147 4379
<< metal4 >>
rect 65 6299 138466 6320
rect 65 4827 138108 6299
rect 65 4654 317 4827
rect 33298 4654 33715 4827
rect 65 4653 33715 4654
rect 137147 4657 138108 4827
rect 138215 4657 138466 6299
rect 137147 4653 138466 4657
rect 65 4635 138466 4653
rect 66 4464 138466 4484
rect 66 4461 33715 4464
rect 66 4288 279 4461
rect 33299 4290 33715 4461
rect 137147 4290 138466 4464
rect 33299 4288 138466 4290
rect 66 2799 138466 4288
<< comment >>
rect 33349 738 33417 817
rect 33827 738 33895 817
rect 33349 580 33895 738
use bias_nstack  bias_nstack_0
array 0 256 -534 0 0 -3895
timestamp 1714090311
transform -1 0 4149 0 -1 1620
box 3258 -2860 3926 1035
use bias_pstack  bias_pstack_0
array 0 256 534 0 0 -4355
timestamp 1714090311
transform 1 0 -1804 0 -1 5026
box 1986 -3967 2714 388
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_3 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform -1 0 147072 0 1 1458
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_5
timestamp 1715205430
transform -1 0 147072 0 1 6342
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_6
timestamp 1715205430
transform -1 0 147072 0 1 4714
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_7
timestamp 1715205430
transform -1 0 147072 0 1 3086
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_8
timestamp 1715205430
transform -1 0 144480 0 1 1458
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_9
timestamp 1715205430
transform -1 0 144480 0 1 4714
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_10
timestamp 1715205430
transform -1 0 144480 0 1 3086
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_11
timestamp 1715205430
transform -1 0 141888 0 1 1458
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_12
timestamp 1715205430
transform -1 0 144480 0 1 6342
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_13
timestamp 1715205430
transform -1 0 141888 0 1 6342
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_14
timestamp 1715205430
transform -1 0 141888 0 -1 3086
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_16
timestamp 1715205430
transform -1 0 141888 0 1 4714
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_17
timestamp 1715205430
transform -1 0 141888 0 1 3086
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_18
timestamp 1715205430
transform -1 0 141888 0 -1 4714
box -66 -43 450 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform -1 0 149280 0 -1 6342
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_1
timestamp 1715205430
transform -1 0 149280 0 -1 3086
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_2
timestamp 1715205430
transform -1 0 149280 0 -1 4714
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_3
timestamp 1715205430
transform -1 0 146688 0 1 1458
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_4
timestamp 1715205430
transform -1 0 149280 0 -1 7970
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_5
timestamp 1715205430
transform -1 0 146688 0 1 6342
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_6
timestamp 1715205430
transform -1 0 146688 0 1 4714
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_7
timestamp 1715205430
transform -1 0 146688 0 1 3086
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_8
timestamp 1715205430
transform -1 0 144096 0 1 1458
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_9
timestamp 1715205430
transform -1 0 144096 0 1 4714
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_10
timestamp 1715205430
transform -1 0 144096 0 1 3086
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_11
timestamp 1715205430
transform -1 0 141504 0 1 1458
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_12
timestamp 1715205430
transform -1 0 144096 0 1 6342
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_13
timestamp 1715205430
transform -1 0 141504 0 1 6342
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_14
timestamp 1715205430
transform -1 0 141504 0 -1 3086
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_16
timestamp 1715205430
transform -1 0 141504 0 1 4714
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_17
timestamp 1715205430
transform -1 0 141504 0 1 3086
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_18
timestamp 1715205430
transform -1 0 141504 0 -1 4714
box -66 -43 162 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform -1 0 147072 0 -1 3086
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_1
timestamp 1715205430
transform -1 0 141888 0 -1 7970
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_5
timestamp 1715205430
transform -1 0 147072 0 -1 7970
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_6
timestamp 1715205430
transform -1 0 147072 0 -1 6342
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_7
timestamp 1715205430
transform -1 0 147072 0 -1 4714
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_8
timestamp 1715205430
transform -1 0 144480 0 -1 4714
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_9
timestamp 1715205430
transform -1 0 144480 0 -1 3086
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_10
timestamp 1715205430
transform -1 0 144480 0 -1 7970
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_11
timestamp 1715205430
transform -1 0 144480 0 -1 6342
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_12
timestamp 1715205430
transform -1 0 141888 0 -1 6342
box -66 -43 546 897
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
array 0 3 -2592 0 3 1628
timestamp 1715205430
transform -1 0 141408 0 1 1458
box -66 -43 2178 1671
<< labels >>
flabel metal3 10199 0 10420 229 0 FreeSans 1600 90 0 0 ena_2000
port 49 nsew
flabel metal3 11094 0 11456 229 0 FreeSans 1600 90 0 0 snk_2000
port 32 nsew
flabel metal2 22467 563 22667 763 0 FreeSans 256 0 0 0 ena
port 11 nsew
flabel metal2 33557 9037 33717 9237 0 FreeSans 256 0 0 0 enb
port 3 nsew
flabel comment 33618 658 33618 658 0 FreeSans 1600 0 0 0 mirror
flabel metal3 41543 9224 41905 9465 0 FreeSans 1600 90 0 0 src_10000_0
port 14 nsew
flabel metal3 40664 9250 40885 9465 0 FreeSans 1600 90 0 0 enb_10000_0
port 13 nsew
flabel metal3 56506 0 56727 229 0 FreeSans 1600 90 0 0 ena_5000_0
port 31 nsew
flabel metal3 57401 0 57763 229 0 FreeSans 1600 90 0 0 snk_5000_0
port 48 nsew
flabel metal3 120882 1 121244 189 0 FreeSans 1600 90 0 0 snk_3700
port 37 nsew
flabel metal3 119987 1 120208 189 0 FreeSans 1600 90 0 0 ena_3700
port 38 nsew
flabel metal3 137060 195 137194 337 0 FreeSans 1600 90 0 0 ena_test1
port 42 nsew
flabel metal3 136670 193 136875 335 0 FreeSans 1600 90 0 0 snk_test1
port 41 nsew
flabel metal3 136664 9225 136907 9466 0 FreeSans 1600 90 0 0 src_test1
port 43 nsew
flabel metal3 137011 9226 137210 9467 0 FreeSans 1600 90 0 0 enb_test1
port 44 nsew
flabel metal3 136322 9225 136543 9465 0 FreeSans 1600 90 0 0 enb_50
port 29 nsew
flabel metal3 135980 9225 136219 9465 0 FreeSans 1600 90 0 0 src_50
port 30 nsew
flabel metal3 135551 9225 135909 9465 0 FreeSans 1600 90 0 0 src_100
port 28 nsew
flabel metal3 135196 9225 135417 9465 0 FreeSans 1600 90 0 0 enb_100
port 27 nsew
flabel metal3 133999 9225 134357 9465 0 FreeSans 1600 90 0 0 src_200_2
port 26 nsew
flabel metal3 133104 9225 133325 9465 0 FreeSans 1600 90 0 0 enb_200_2
port 25 nsew
flabel metal3 131907 9225 132265 9465 0 FreeSans 1600 90 0 0 src_200_1
port 24 nsew
flabel metal3 131012 9225 131233 9465 0 FreeSans 1600 90 0 0 enb_200_1
port 23 nsew
flabel metal3 129815 9225 130173 9465 0 FreeSans 1600 90 0 0 src_200_0
port 22 nsew
flabel metal3 128920 9225 129141 9465 0 FreeSans 1600 90 0 0 enb_200_0
port 21 nsew
flabel metal3 126645 9225 127003 9465 0 FreeSans 1600 90 0 0 src_400
port 20 nsew
flabel metal3 125750 9225 125971 9465 0 FreeSans 1600 90 0 0 enb_400
port 19 nsew
flabel metal3 121385 9224 121747 9465 0 FreeSans 1600 90 0 0 src_600
port 18 nsew
flabel metal3 120490 9225 120711 9466 0 FreeSans 1600 90 0 0 enb_600
port 17 nsew
flabel metal3 64774 1 65136 230 0 FreeSans 1600 90 0 0 snk_5000_2
port 36 nsew
flabel metal3 63879 1 64100 230 0 FreeSans 1600 90 0 0 ena_5000_2
port 35 nsew
flabel metal3 54217 9224 54579 9465 0 FreeSans 1600 90 0 0 src_10000_1
port 15 nsew
flabel metal3 53322 9224 53543 9465 0 FreeSans 1600 90 0 0 enb_10000_1
port 16 nsew
flabel metal4 65 4635 298 6320 0 FreeSans 1600 90 0 0 avdd
port 47 nsew
flabel metal4 66 2799 299 4484 0 FreeSans 1600 90 0 0 avss
port 12 nsew
<< end >>
