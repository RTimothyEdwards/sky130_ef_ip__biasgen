magic
tech sky130A
magscale 1 2
timestamp 1716925149
<< pwell >>
rect -715 -458 715 458
<< mvnmos >>
rect -487 -200 -287 200
rect -229 -200 -29 200
rect 29 -200 229 200
rect 287 -200 487 200
<< mvndiff >>
rect -545 188 -487 200
rect -545 -188 -533 188
rect -499 -188 -487 188
rect -545 -200 -487 -188
rect -287 188 -229 200
rect -287 -188 -275 188
rect -241 -188 -229 188
rect -287 -200 -229 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 229 188 287 200
rect 229 -188 241 188
rect 275 -188 287 188
rect 229 -200 287 -188
rect 487 188 545 200
rect 487 -188 499 188
rect 533 -188 545 188
rect 487 -200 545 -188
<< mvndiffc >>
rect -533 -188 -499 188
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
rect 499 -188 533 188
<< mvpsubdiff >>
rect -679 410 679 422
rect -679 376 -571 410
rect 571 376 679 410
rect -679 364 679 376
rect -679 314 -621 364
rect -679 -314 -667 314
rect -633 -314 -621 314
rect 621 314 679 364
rect -679 -364 -621 -314
rect 621 -314 633 314
rect 667 -314 679 314
rect 621 -364 679 -314
rect -679 -376 679 -364
rect -679 -410 -571 -376
rect 571 -410 679 -376
rect -679 -422 679 -410
<< mvpsubdiffcont >>
rect -571 376 571 410
rect -667 -314 -633 314
rect 633 -314 667 314
rect -571 -410 571 -376
<< poly >>
rect -487 272 -287 288
rect -487 238 -471 272
rect -303 238 -287 272
rect -487 200 -287 238
rect -229 272 -29 288
rect -229 238 -213 272
rect -45 238 -29 272
rect -229 200 -29 238
rect 29 272 229 288
rect 29 238 45 272
rect 213 238 229 272
rect 29 200 229 238
rect 287 272 487 288
rect 287 238 303 272
rect 471 238 487 272
rect 287 200 487 238
rect -487 -238 -287 -200
rect -487 -272 -471 -238
rect -303 -272 -287 -238
rect -487 -288 -287 -272
rect -229 -238 -29 -200
rect -229 -272 -213 -238
rect -45 -272 -29 -238
rect -229 -288 -29 -272
rect 29 -238 229 -200
rect 29 -272 45 -238
rect 213 -272 229 -238
rect 29 -288 229 -272
rect 287 -238 487 -200
rect 287 -272 303 -238
rect 471 -272 487 -238
rect 287 -288 487 -272
<< polycont >>
rect -471 238 -303 272
rect -213 238 -45 272
rect 45 238 213 272
rect 303 238 471 272
rect -471 -272 -303 -238
rect -213 -272 -45 -238
rect 45 -272 213 -238
rect 303 -272 471 -238
<< locali >>
rect -667 376 -571 410
rect 571 376 667 410
rect -667 314 -633 376
rect 633 314 667 376
rect -487 238 -471 272
rect -303 238 -287 272
rect -229 238 -213 272
rect -45 238 -29 272
rect 29 238 45 272
rect 213 238 229 272
rect 287 238 303 272
rect 471 238 487 272
rect -533 188 -499 204
rect -533 -204 -499 -188
rect -275 188 -241 204
rect -275 -204 -241 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 241 188 275 204
rect 241 -204 275 -188
rect 499 188 533 204
rect 499 -204 533 -188
rect -487 -272 -471 -238
rect -303 -272 -287 -238
rect -229 -272 -213 -238
rect -45 -272 -29 -238
rect 29 -272 45 -238
rect 213 -272 229 -238
rect 287 -272 303 -238
rect 471 -272 487 -238
rect -667 -376 -633 -314
rect 633 -376 667 -314
rect -667 -410 -571 -376
rect 571 -410 667 -376
<< viali >>
rect -450 238 -324 272
rect -192 238 -66 272
rect 66 238 192 272
rect 324 238 450 272
rect -533 -188 -499 188
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
rect 499 -188 533 188
rect -450 -272 -324 -238
rect -192 -272 -66 -238
rect 66 -272 192 -238
rect 324 -272 450 -238
<< metal1 >>
rect -462 272 -312 278
rect -462 238 -450 272
rect -324 238 -312 272
rect -462 232 -312 238
rect -204 272 -54 278
rect -204 238 -192 272
rect -66 238 -54 272
rect -204 232 -54 238
rect 54 272 204 278
rect 54 238 66 272
rect 192 238 204 272
rect 54 232 204 238
rect 312 272 462 278
rect 312 238 324 272
rect 450 238 462 272
rect 312 232 462 238
rect -539 188 -493 200
rect -539 -188 -533 188
rect -499 -188 -493 188
rect -539 -200 -493 -188
rect -281 188 -235 200
rect -281 -188 -275 188
rect -241 -188 -235 188
rect -281 -200 -235 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 235 188 281 200
rect 235 -188 241 188
rect 275 -188 281 188
rect 235 -200 281 -188
rect 493 188 539 200
rect 493 -188 499 188
rect 533 -188 539 188
rect 493 -200 539 -188
rect -462 -238 -312 -232
rect -462 -272 -450 -238
rect -324 -272 -312 -238
rect -462 -278 -312 -272
rect -204 -238 -54 -232
rect -204 -272 -192 -238
rect -66 -272 -54 -238
rect -204 -278 -54 -272
rect 54 -238 204 -232
rect 54 -272 66 -238
rect 192 -272 204 -238
rect 54 -278 204 -272
rect 312 -238 462 -232
rect 312 -272 324 -238
rect 450 -272 462 -238
rect 312 -278 462 -272
<< properties >>
string FIXED_BBOX -650 -393 650 393
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2 l 1 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 75 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
