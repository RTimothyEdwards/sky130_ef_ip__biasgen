magic
tech sky130A
magscale 1 2
timestamp 1716925149
<< error_s >>
rect 5281 5205 8276 5386
rect 5281 5100 5736 5205
rect 6710 5100 8276 5205
rect 5281 2686 5567 5100
rect 7990 2686 8276 5100
rect 5281 2400 8276 2686
<< dnwell >>
rect 5361 2480 8196 5306
<< viali >>
rect 5921 5099 6523 5143
rect 5641 3169 6784 3223
<< metal1 >>
rect 5901 5150 6547 5161
rect 5901 5093 5910 5150
rect 6536 5093 6547 5150
rect 5901 5083 6547 5093
rect 5911 4465 5951 4895
rect 6016 4465 6044 4988
rect 6074 4893 6372 4910
rect 6074 4809 6092 4893
rect 6359 4809 6372 4893
rect 6074 4793 6372 4809
rect 6402 4465 6430 4986
rect 5911 4428 6015 4465
rect 6016 4428 6448 4465
rect 5557 4068 5590 4347
rect 5911 4171 5951 4428
rect 6489 4175 6529 4905
rect 5911 4131 5975 4171
rect 5557 4035 5890 4068
rect 5615 3781 5827 3794
rect 5615 3686 5632 3781
rect 5809 3686 5827 3781
rect 5615 3673 5827 3686
rect 5857 3345 5890 4035
rect 5935 3576 5975 4131
rect 6452 4135 6529 4175
rect 5901 3320 6012 3366
rect 6033 3341 6066 3858
rect 6099 3777 6321 3792
rect 6099 3682 6115 3777
rect 6302 3682 6321 3777
rect 6099 3671 6321 3682
rect 6367 3337 6400 3854
rect 6452 3578 6492 4135
rect 6789 4066 6822 4339
rect 6535 4033 6822 4066
rect 6416 3320 6527 3366
rect 6535 3339 6568 4033
rect 6596 3780 6798 3796
rect 6596 3685 6613 3780
rect 6780 3685 6798 3780
rect 6596 3675 6798 3685
rect 6958 3506 7183 3524
rect 6958 3416 6974 3506
rect 7163 3416 7183 3506
rect 6958 3401 7183 3416
rect 5627 3223 6797 3233
rect 5627 3169 5641 3223
rect 6784 3169 6797 3223
rect 5627 3158 6797 3169
rect 7212 3038 7245 3852
rect 7291 3557 7606 3648
rect 7187 3030 7276 3038
rect 7187 2808 7195 3030
rect 7267 2808 7276 3030
rect 7187 2800 7276 2808
rect 7655 2708 7688 3851
rect 7716 3778 7946 3794
rect 7716 3690 7732 3778
rect 7929 3690 7946 3778
rect 7716 3674 7946 3690
rect 7526 2699 7692 2708
rect 7526 2647 7534 2699
rect 7683 2647 7692 2699
rect 7526 2639 7692 2647
<< via1 >>
rect 5910 5143 6536 5150
rect 5910 5099 5921 5143
rect 5921 5099 6523 5143
rect 6523 5099 6536 5143
rect 5910 5093 6536 5099
rect 6092 4809 6359 4893
rect 5632 3686 5809 3781
rect 6115 3682 6302 3777
rect 6613 3685 6780 3780
rect 6974 3416 7163 3506
rect 5641 3169 6784 3223
rect 7195 2808 7267 3030
rect 7732 3690 7929 3778
rect 7534 2647 7683 2699
<< metal2 >>
rect 5443 5156 7868 5172
rect 5443 5150 7112 5156
rect 5443 5093 5910 5150
rect 6536 5093 7112 5150
rect 5443 4893 7112 5093
rect 5443 4809 6092 4893
rect 6359 4809 7112 4893
rect 5443 4802 7112 4809
rect 7851 4802 7868 5156
rect 5443 4785 7868 4802
rect 5530 3781 7960 3959
rect 5530 3686 5632 3781
rect 5809 3780 7960 3781
rect 5809 3777 6613 3780
rect 5809 3686 6115 3777
rect 5530 3682 6115 3686
rect 6302 3685 6613 3777
rect 6780 3778 7960 3780
rect 6780 3690 7732 3778
rect 7929 3690 7960 3778
rect 6780 3685 7960 3690
rect 6302 3682 7960 3685
rect 5530 3671 7960 3682
rect 5476 3506 7956 3521
rect 5476 3416 6974 3506
rect 7163 3501 7956 3506
rect 7163 3416 7204 3501
rect 5476 3223 7204 3416
rect 5476 3169 5641 3223
rect 6784 3169 7204 3223
rect 5476 3165 7204 3169
rect 7930 3165 7956 3501
rect 5476 3146 7956 3165
rect 5480 3030 8196 3038
rect 5480 2808 7195 3030
rect 7267 2808 8196 3030
rect 5480 2800 8196 2808
rect 7526 2699 7692 2708
rect 7526 2684 7534 2699
rect 5495 2647 7534 2684
rect 7683 2647 7692 2699
rect 5495 2646 7692 2647
rect 7526 2639 7692 2646
<< via2 >>
rect 7112 4802 7851 5156
rect 7204 3165 7930 3501
<< metal3 >>
rect 7094 5156 7868 5172
rect 7094 4802 7112 5156
rect 7851 4802 7868 5156
rect 7094 4784 7868 4802
rect 7179 3501 7955 3522
rect 7179 3165 7204 3501
rect 7930 3165 7955 3501
rect 7179 3147 7955 3165
use sky130_fd_pr__nfet_05v0_nvt_F3TL5C  sky130_fd_pr__nfet_05v0_nvt_F3TL5C_0 paramcells
timestamp 1716925149
transform 1 0 7733 0 -1 3598
box -328 -458 328 458
use sky130_fd_pr__nfet_g5v0d10v5_56WC32  sky130_fd_pr__nfet_g5v0d10v5_56WC32_0 paramcells
timestamp 1716925149
transform 1 0 7167 0 -1 3598
box -368 -458 368 458
use sky130_fd_pr__nfet_g5v0d10v5_V5WCXY  sky130_fd_pr__nfet_g5v0d10v5_V5WCXY_0 paramcells
timestamp 1716925149
transform 1 0 6214 0 -1 3598
box -715 -458 715 458
use sky130_fd_pr__pfet_g5v0d10v5_QSDYAY  sky130_fd_pr__pfet_g5v0d10v5_QSDYAY_0 paramcells
timestamp 1716912327
transform 1 0 6223 0 -1 4708
box -487 -497 487 497
<< labels >>
flabel metal2 5443 4785 5725 5073 0 FreeSans 1600 0 0 0 avdd
port 1 nsew
flabel metal2 5480 2800 5707 3038 0 FreeSans 800 0 0 0 nbias
port 2 nsew
flabel metal2 5495 2646 5784 2684 0 FreeSans 320 0 0 0 ena
port 3 nsew
flabel metal2 5476 3233 5784 3521 0 FreeSans 1600 0 0 0 avss
port 4 nsew
flabel metal1 5557 4211 5590 4347 0 FreeSans 320 90 0 0 inp
port 5 nsew
flabel metal1 6789 4203 6822 4339 0 FreeSans 320 90 0 0 inn
port 6 nsew
<< end >>
