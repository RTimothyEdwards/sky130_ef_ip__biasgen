magic
tech sky130A
magscale 1 2
timestamp 1716925370
<< error_s >>
rect 45862 8386 45886 8410
rect 45886 8352 45910 8386
rect 45862 8328 45886 8352
rect 45886 8233 45952 8262
rect 45886 8200 45966 8233
rect 45862 8196 45966 8200
rect 45820 8153 45966 8196
rect 44986 7494 45966 8153
rect 20242 6143 20244 7195
rect 44986 7047 45886 7494
rect 20036 5937 20450 6143
rect 20036 5935 21502 5937
rect 20036 5729 20450 5935
rect 45885 4320 45886 4409
rect 45881 4292 45886 4320
rect 45905 4292 45966 7494
rect 44986 3392 45966 4292
rect 45680 507 45966 3392
rect 45886 336 45966 507
rect 45862 332 45966 336
rect 45820 258 45966 332
rect 45862 254 45966 258
rect 45886 221 45966 254
rect 45886 192 45952 221
rect 45880 104 45886 105
rect 45862 80 45886 104
rect 45880 61 45910 80
rect 45886 46 45910 61
rect 45862 22 45886 46
<< dnwell >>
rect 5006 5937 45886 8153
rect 5006 5935 20242 5937
rect 20244 5935 45886 5937
rect 5006 301 45886 5935
<< nwell >>
rect 4897 7947 45886 8262
rect 4897 507 5212 7947
rect 4897 192 45886 507
<< pwell >>
rect 19789 766 19859 1198
rect 35342 507 35430 529
<< mvpsubdiff >>
rect 4777 8352 4837 8386
rect 4777 8326 4811 8352
rect 1075 7702 1135 7736
rect 4170 7702 4230 7736
rect 1075 7676 1109 7702
rect 1075 682 1109 708
rect 4196 7676 4230 7702
rect 4196 682 4230 708
rect 1075 648 1135 682
rect 4170 648 4230 682
rect 4777 80 4811 106
rect 4777 46 4837 80
<< mvnsubdiff >>
rect 4963 8176 45886 8196
rect 4963 8142 5043 8176
rect 4963 8122 45886 8142
rect 4963 8116 5037 8122
rect 4963 338 4983 8116
rect 5017 338 5037 8116
rect 4963 332 5037 338
rect 4963 312 45886 332
rect 4963 278 5043 312
rect 4963 258 45886 278
<< mvpsubdiffcont >>
rect 4837 8352 45886 8386
rect 1135 7702 4170 7736
rect 1075 708 1109 7676
rect 4196 708 4230 7676
rect 1135 648 4170 682
rect 4777 106 4811 8326
rect 4837 46 45886 80
<< mvnsubdiffcont >>
rect 5043 8142 45886 8176
rect 4983 338 5017 8116
rect 5043 278 45886 312
<< locali >>
rect 4777 8352 4837 8386
rect 4777 8326 45886 8352
rect 1072 7736 4777 7837
rect 1072 7702 1135 7736
rect 4170 7713 4777 7736
rect 4170 7702 4341 7713
rect 1072 7676 1209 7702
rect 1072 708 1075 7676
rect 1109 708 1209 7676
rect 4196 7676 4341 7702
rect 3464 7097 3511 7163
rect 1707 6273 1873 6285
rect 1707 6164 1720 6273
rect 1857 6164 1873 6273
rect 1707 6151 1873 6164
rect 1707 4645 1873 4657
rect 1707 4536 1720 4645
rect 1857 4536 1873 4645
rect 1707 4523 1873 4536
rect 3464 3841 3511 3907
rect 1707 3017 1873 3029
rect 1707 2908 1720 3017
rect 1857 2908 1873 3017
rect 1707 2895 1873 2908
rect 1707 1389 1873 1401
rect 1707 1280 1720 1389
rect 1857 1280 1873 1389
rect 1707 1267 1873 1280
rect 1072 682 1209 708
rect 4230 708 4341 7676
rect 4196 682 4341 708
rect 4811 8253 45886 8326
rect 4811 2306 4879 8253
rect 1072 648 1135 682
rect 4170 648 4777 682
rect 1072 558 4777 648
rect 4852 224 4879 2306
rect 4983 8142 5043 8176
rect 4983 8116 45886 8142
rect 5017 7957 45886 8116
rect 5017 7498 5151 7957
rect 5136 7294 5151 7498
rect 5017 491 5151 7294
rect 5017 338 45886 491
rect 4983 312 45886 338
rect 4983 278 5043 312
rect 4811 192 4879 224
rect 4811 106 45886 192
rect 4777 105 45886 106
rect 4777 61 4804 105
rect 4777 46 4837 61
<< viali >>
rect 3782 7073 3848 7300
rect 3398 6825 3464 7052
rect 1720 6164 1857 6273
rect 3398 5197 3464 5424
rect 1720 4536 1857 4645
rect 3782 3817 3848 4044
rect 1720 2908 1857 3017
rect 3398 1941 3464 2168
rect 1720 1280 1857 1389
rect 4803 224 4811 2306
rect 4811 224 4852 2306
rect 4999 7294 5017 7498
rect 5017 7294 5136 7498
rect 4804 80 45886 105
rect 4804 61 4837 80
rect 4837 61 45886 80
<< metal1 >>
rect 19595 8229 19795 8502
rect 19859 7753 33103 7764
rect 19859 7701 19892 7753
rect 33067 7701 33103 7753
rect 19859 7689 33103 7701
rect 4982 7498 5151 7512
rect 3775 7300 3856 7317
rect 3775 7073 3782 7300
rect 3848 7175 3856 7300
rect 4982 7294 4999 7498
rect 5136 7294 5151 7498
rect 4982 7278 5151 7294
rect 3848 7112 4568 7175
rect 3848 7073 3856 7112
rect 3391 7052 3472 7069
rect 3775 7060 3856 7073
rect 3391 6825 3398 7052
rect 3464 6938 3472 7052
rect 3464 6880 4574 6938
rect 3464 6825 3472 6880
rect 3391 6812 3472 6825
rect 1707 6273 1873 6285
rect 1707 6253 1720 6273
rect 1072 6185 1720 6253
rect 1707 6164 1720 6185
rect 1857 6164 1873 6273
rect 1707 6151 1873 6164
rect 3391 5424 3472 5441
rect 3391 5197 3398 5424
rect 3464 5310 3472 5424
rect 3464 5252 4574 5310
rect 3464 5197 3472 5252
rect 3391 5184 3472 5197
rect 1707 4645 1873 4657
rect 1707 4625 1720 4645
rect 1072 4557 1720 4625
rect 1707 4536 1720 4557
rect 1857 4536 1873 4645
rect 1707 4523 1873 4536
rect 3775 4044 3856 4061
rect 3775 3817 3782 4044
rect 3848 3921 3856 4044
rect 3848 3864 4507 3921
rect 3848 3817 3856 3864
rect 3775 3804 3856 3817
rect 1707 3017 1873 3029
rect 1707 2997 1720 3017
rect 1072 2929 1720 2997
rect 1707 2908 1720 2929
rect 1857 2908 1873 3017
rect 1707 2895 1873 2908
rect 4777 2306 4879 2345
rect 3391 2168 3472 2185
rect 4777 2181 4803 2306
rect 3391 1941 3398 2168
rect 3464 2054 3472 2168
rect 3464 1996 4574 2054
rect 3464 1941 3472 1996
rect 3391 1928 3472 1941
rect 1707 1389 1873 1401
rect 1707 1369 1720 1389
rect 1072 1301 1720 1369
rect 1707 1280 1720 1301
rect 1857 1280 1873 1389
rect 1707 1267 1873 1280
rect 4775 622 4803 2181
rect 4777 224 4803 622
rect 4852 2181 4879 2306
rect 4852 2161 5211 2181
rect 4852 641 5042 2161
rect 5198 641 5211 2161
rect 4852 622 5211 641
rect 19541 1066 19593 7598
rect 19653 7166 19859 7598
rect 19955 7166 20191 7598
rect 20287 7166 20523 7598
rect 20619 7166 20855 7598
rect 20951 7166 21187 7598
rect 21283 7166 21519 7598
rect 21615 7166 21851 7598
rect 21947 7166 22183 7598
rect 22279 7166 22515 7598
rect 22611 7166 22847 7598
rect 22943 7166 23179 7598
rect 23275 7166 23511 7598
rect 23607 7166 23843 7598
rect 23939 7166 24175 7598
rect 24271 7166 24507 7598
rect 24603 7166 24839 7598
rect 24935 7166 25171 7598
rect 25267 7166 25503 7598
rect 25599 7166 25835 7598
rect 25931 7166 26167 7598
rect 26263 7166 26499 7598
rect 26595 7166 26831 7598
rect 26927 7166 27163 7598
rect 27259 7166 27495 7598
rect 27591 7166 27827 7598
rect 19541 630 19593 828
rect 19653 1066 19705 7004
rect 27923 6512 28159 7598
rect 28255 7166 28491 7598
rect 28587 7166 28823 7598
rect 28919 7166 29155 7598
rect 29251 7166 29487 7598
rect 29583 7166 29819 7598
rect 29915 7166 30151 7598
rect 30247 7166 30483 7598
rect 30579 7166 30815 7598
rect 30911 7166 31147 7598
rect 31243 7166 31479 7598
rect 31575 7166 31811 7598
rect 31907 7166 32143 7598
rect 32239 7166 32475 7598
rect 32571 7166 32807 7598
rect 32902 7306 33103 7598
rect 32902 7166 33350 7306
rect 27923 6263 28159 6278
rect 33063 4062 33115 4076
rect 33063 3810 33115 3824
rect 33210 2196 33350 7166
rect 33210 1673 33350 1710
rect 19653 630 19705 828
rect 19789 766 20025 1198
rect 20121 766 20357 1198
rect 20453 766 20689 1198
rect 20785 766 21021 1198
rect 21117 766 21353 1198
rect 21449 766 21685 1198
rect 21781 766 22017 1198
rect 22113 766 22349 1198
rect 22445 766 22681 1198
rect 22777 766 23013 1198
rect 23109 766 23345 1198
rect 23441 766 23677 1198
rect 23773 766 24009 1198
rect 24105 766 24341 1198
rect 24437 766 24673 1198
rect 24769 766 25005 1198
rect 25101 766 25337 1198
rect 25433 766 25669 1198
rect 25765 766 26001 1198
rect 26097 766 26333 1198
rect 26429 766 26665 1198
rect 26761 766 26997 1198
rect 27093 766 27329 1198
rect 27425 766 27661 1198
rect 27757 766 27993 1198
rect 28089 766 28325 1198
rect 28421 766 28657 1198
rect 28753 766 28989 1198
rect 29085 766 29321 1198
rect 29417 766 29653 1198
rect 29749 766 29985 1198
rect 30081 766 30317 1198
rect 30413 766 30649 1198
rect 30745 766 30981 1198
rect 31077 766 31313 1198
rect 31409 766 31645 1198
rect 31741 766 31977 1198
rect 32073 766 32309 1198
rect 32405 766 32641 1198
rect 32737 766 32973 1198
rect 33063 630 33109 1360
rect 4852 224 4879 622
rect 4777 124 4879 224
rect 4777 105 45886 124
rect 4777 61 4804 105
rect 4777 46 45886 61
<< via1 >>
rect 19892 7701 33067 7753
rect 4999 7294 5136 7498
rect 5042 641 5198 2161
rect 19541 828 19593 1066
rect 27923 6278 28159 6512
rect 33063 3824 33115 4062
rect 33210 1710 33350 2196
rect 19653 828 19705 1066
<< metal2 >>
rect 33578 8317 33721 8549
rect 33927 8317 34186 8549
rect 34631 8317 45886 8549
rect 33764 8010 34057 8242
rect 34263 8010 34362 8242
rect 34631 8010 45886 8242
rect 5108 7753 33185 7847
rect 5108 7701 19892 7753
rect 33067 7701 33185 7753
rect 5108 7609 33185 7701
rect 33426 7609 45886 7847
rect 4982 7498 33435 7512
rect 4982 7294 4999 7498
rect 5136 7294 33435 7498
rect 4982 7278 33435 7294
rect 19586 6278 27923 6512
rect 28159 6278 45886 6512
rect 33202 6277 33433 6278
rect 5477 5274 45886 5508
rect 33053 3824 33063 4062
rect 33115 3824 33186 4062
rect 33427 4043 34526 4062
rect 33427 3959 33565 4043
rect 33427 3824 34526 3959
rect 8196 2800 45886 3038
rect 4775 2161 5211 2181
rect 4775 641 5042 2161
rect 5198 1066 5211 2161
rect 33198 1710 33210 2196
rect 33350 2054 33361 2196
rect 33350 1816 45886 2054
rect 33350 1710 33361 1816
rect 33198 1709 33361 1710
rect 5198 828 19541 1066
rect 19593 828 19653 1066
rect 19705 828 33186 1066
rect 33427 828 45886 1066
rect 5198 641 5211 828
rect 4775 622 5211 641
rect 33157 431 33186 619
rect 33312 431 34367 619
rect 34435 431 45886 619
rect 33597 175 33783 363
rect 33983 175 34207 363
rect 34654 175 44951 363
rect 45301 175 45653 363
<< via2 >>
rect 33721 8317 33927 8549
rect 34057 8010 34263 8242
rect 33185 7609 33426 7847
rect 33564 4236 45886 4320
rect 33186 3824 33427 4062
rect 33565 3959 45886 4043
rect 5042 641 5198 2161
rect 33186 828 33427 1066
rect 33186 431 33312 619
rect 33783 175 33983 363
<< metal3 >>
rect 33709 8549 33938 8863
rect 33709 8317 33721 8549
rect 33927 8317 33938 8549
rect 33709 8304 33938 8317
rect 34045 8242 34274 8863
rect 34045 8010 34057 8242
rect 34263 8010 34274 8242
rect 34045 7994 34274 8010
rect 33175 7847 33437 7875
rect 33175 7609 33185 7847
rect 33426 7609 33437 7847
rect 33175 4062 33437 7609
rect 33539 4409 45886 4454
rect 33539 4236 33564 4409
rect 33539 4220 45886 4236
rect 33175 3824 33186 4062
rect 33427 4043 45886 4062
rect 33427 3870 33521 4043
rect 33427 3824 45886 3870
rect 4775 2161 5211 2181
rect 4775 641 5042 2161
rect 5198 641 5211 2161
rect 33175 1066 33437 3824
rect 33175 828 33186 1066
rect 33427 828 33437 1066
rect 33175 794 33437 828
rect 4775 622 5211 641
rect 33179 619 33319 627
rect 33179 431 33186 619
rect 33312 431 33319 619
rect 33179 159 33319 431
rect 33776 363 33991 385
rect 33776 175 33783 363
rect 33983 175 33991 363
rect 33776 0 33991 175
<< via3 >>
rect 7112 4802 7851 5156
rect 33564 4320 45886 4409
rect 33564 4236 45886 4320
rect 33521 3959 33565 4043
rect 33565 3959 45886 4043
rect 33521 3870 45886 3959
rect 7204 3165 7930 3501
rect 5042 641 5198 2161
<< metal4 >>
rect 4770 5156 45886 5902
rect 4770 4802 7112 5156
rect 7851 4802 45886 5156
rect 4770 4409 45886 4802
rect 4770 4236 33564 4409
rect 4770 4217 45886 4236
rect 4777 4043 45886 4066
rect 4777 3870 33521 4043
rect 4777 3501 45886 3870
rect 4777 3165 7204 3501
rect 7930 3165 45886 3501
rect 4777 2381 45886 3165
rect 4775 2161 5211 2182
rect 4775 641 5042 2161
rect 5198 641 5211 2161
rect 4775 622 5211 641
use bias_amp  bias_amp_0
timestamp 1716925149
transform 1 0 0 0 1 0
box 5281 2400 8276 5386
use bias_nstack  bias_nstack_0
array 0 22 -534 0 0 -3895
timestamp 1714090311
transform -1 0 37396 0 -1 1202
box 3258 -2860 3926 1035
use bias_pstack  bias_pstack_0
array 0 22 534 0 0 -4355
timestamp 1714090311
transform 1 0 31443 0 -1 4608
box 1986 -3967 2714 388
use sky130_fd_pr__cap_mim_m3_1_MQZGVK  sky130_fd_pr__cap_mim_m3_1_MQZGVK_0 paramcells
timestamp 1716925149
transform 0 1 8149 1 0 6878
box -686 -2640 686 2640
use sky130_fd_pr__cap_mim_m3_1_MQZGVK  sky130_fd_pr__cap_mim_m3_1_MQZGVK_1
timestamp 1716925149
transform 0 1 8170 -1 0 1389
box -686 -2640 686 2640
use sky130_fd_pr__res_high_po_0p35_L4QTBM  sky130_fd_pr__res_high_po_0p35_L4QTBM_0 paramcells
timestamp 1716925149
transform 1 0 13944 0 1 4182
box -5679 -3582 5679 3582
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform 1 0 3486 0 1 4217
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_1
timestamp 1715205430
transform 1 0 3486 0 1 961
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_2
timestamp 1715205430
transform 1 0 3486 0 1 2589
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_3
timestamp 1715205430
transform 1 0 3486 0 -1 5845
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_4
timestamp 1715205430
transform 1 0 3486 0 1 5845
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_11
timestamp 1715205430
transform 1 0 3486 0 -1 2589
box -66 -43 450 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform 1 0 3870 0 1 4217
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_1
timestamp 1715205430
transform 1 0 3870 0 -1 2589
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_2
timestamp 1715205430
transform 1 0 3870 0 1 2589
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_3
timestamp 1715205430
transform 1 0 3870 0 -1 5845
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_4
timestamp 1715205430
transform 1 0 3870 0 1 5845
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_11
timestamp 1715205430
transform 1 0 3870 0 1 961
box -66 -43 162 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_2 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform 1 0 3486 0 -1 4217
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_4
timestamp 1715205430
transform 1 0 3486 0 -1 7473
box -66 -43 546 897
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
array 0 0 2592 0 3 1628
timestamp 1715205430
transform 1 0 1374 0 1 961
box -66 -43 2178 1671
use sky130_fd_pr__res_high_po_0p35_P35QVK  XR2 paramcells
timestamp 1713888873
transform 1 0 26381 0 1 4182
box -6758 -3582 6758 3582
<< labels >>
flabel metal3 33179 159 33319 296 0 FreeSans 1600 90 0 0 ena_test0
port 39 nsew
flabel metal3 33776 0 33991 153 0 FreeSans 1600 90 0 0 snk_test0
port 40 nsew
flabel metal3 33709 8630 33938 8863 0 FreeSans 1600 90 0 0 src_test0
port 45 nsew
flabel metal3 34045 8630 34274 8863 0 FreeSans 1600 90 0 0 enb_test0
port 46 nsew
flabel metal4 4770 4217 5003 5902 0 FreeSans 1600 90 0 0 avdd
port 47 nsew
flabel metal4 4777 2381 5010 4066 0 FreeSans 1600 90 0 0 avss
port 12 nsew
flabel metal4 4775 622 5042 2182 0 FreeSans 1600 90 0 0 vsub
port 50 nsew
flabel metal1 19595 8302 19795 8502 0 FreeSans 256 90 0 0 ref_in
port 1 nsew
flabel metal1 1072 6185 1472 6253 0 FreeSans 480 0 0 0 ref_sel_vbg
port 52 nsew
flabel metal1 1072 4557 1472 4625 0 FreeSans 480 0 0 0 ena
port 53 nsew
flabel metal1 1072 2929 1472 2997 0 FreeSans 480 0 0 0 ena_src_test0
port 54 nsew
flabel metal1 1072 1301 1472 1369 0 FreeSans 480 0 0 0 ena_snk_test0
port 55 nsew
flabel metal1 4150 3892 4150 3892 0 FreeSans 480 0 0 0 enb_test0_3v3
flabel metal1 4127 5281 4127 5281 0 FreeSans 480 0 0 0 ena_3v3
flabel metal1 4052 2022 4052 2022 0 FreeSans 480 0 0 0 ena_test0_3v3
flabel metal1 4118 6906 4118 6906 0 FreeSans 480 0 0 0 ena_vbg_3v3
flabel metal1 4133 7133 4133 7133 0 FreeSans 480 0 0 0 enb_vbg_3v3
<< end >>
