magic
tech sky130A
magscale 1 2
timestamp 1717075507
<< metal1 >>
rect 5441 8326 5562 8557
rect 1072 6185 1472 6253
rect 1072 4557 1472 4625
rect 1072 2929 1472 2997
rect 1072 1301 1472 1369
<< metal2 >>
rect 4682 2646 5538 2684
use bias_generator_be  bias_generator_be_0
timestamp 1717075507
transform 1 0 45529 0 1 -418
box -24 0 149476 9467
use bias_generator_fe  bias_generator_fe_0
timestamp 1717075507
transform 1 0 0 0 1 0
box 1072 0 45976 8863
<< labels >>
flabel metal1 1072 6185 1472 6253 0 FreeSans 480 0 0 0 ref_sel_vbg
port 52 nsew
flabel metal1 1072 4557 1472 4625 0 FreeSans 480 0 0 0 ena
port 53 nsew
flabel metal1 1072 2929 1472 2997 0 FreeSans 480 0 0 0 ena_src_test0
port 54 nsew
flabel metal1 1072 1301 1472 1369 0 FreeSans 480 0 0 0 ena_snk_test0
port 55 nsew
flabel metal1 5441 8326 5562 8557 0 FreeSans 1600 90 0 0 vbg
port 56 nsew
<< end >>
